rommem[0] = 33'h0C2FB1878;
rommem[1] = 33'h0DFFFA230;
rommem[2] = 33'h0FA33A09A;
rommem[3] = 33'h0290000B9;
rommem[4] = 33'h00CF000FF;
rommem[5] = 33'h09FF00009;
rommem[6] = 33'h0E8F10040;
rommem[7] = 33'h1EC80C8E8;
rommem[8] = 33'h1FFA9DE80;
rommem[9] = 33'h1E0308DFF;
rommem[10] = 33'h126642464;
rommem[11] = 33'h1850014A9;
rommem[12] = 33'h000F1A92C;
rommem[13] = 33'h110642E85;
rommem[14] = 33'h1F0A91464;
rommem[15] = 33'h1A9128500;
rommem[16] = 33'h1168500F1;
rommem[17] = 33'h1850014A9;
rommem[18] = 33'h0A91A6414;
rommem[19] = 33'h13085001D;
rommem[20] = 33'h0850038A9;
rommem[21] = 33'h10099A934;
rommem[22] = 33'h0A903008D;
rommem[23] = 33'h1028D00F0;
rommem[24] = 33'h0A93E6403;
rommem[25] = 33'h13C85FA33;
rommem[26] = 33'h0CBF2AE20;
rommem[27] = 33'h1AD20E208;
rommem[28] = 33'h129AAF06F;
rommem[29] = 33'h18A1BD001;
rommem[30] = 33'h103D00229;
rommem[31] = 33'h08DEC8028;
rommem[32] = 33'h1E628F07E;
rommem[33] = 33'h1E602D024;
rommem[34] = 33'h00020A926;
rommem[35] = 33'h11A641485;
rommem[36] = 33'h0908DD980;
rommem[37] = 33'h1004C28F0;
rommem[38] = 33'h000FF29F8;
rommem[39] = 33'h137302824;
rommem[40] = 33'h1F00008C9;
rommem[41] = 33'h10091C935;
rommem[42] = 33'h093C933F0;
rommem[43] = 33'h1C931F000;
rommem[44] = 33'h12FF00090;
rommem[45] = 33'h1F00092C9;
rommem[46] = 33'h00099C92D;
rommem[47] = 33'h10DC92BF0;
rommem[48] = 33'h1C957F000;
rommem[49] = 33'h157F0000A;
rommem[50] = 33'h1F00094C9;
rommem[51] = 33'h1001BC91F;
rommem[52] = 33'h028641DD0;
rommem[53] = 33'h0826028C6;
rommem[54] = 33'h000820053;
rommem[55] = 33'h1014A8201;
rommem[56] = 33'h082015282;
rommem[57] = 33'h15A820156;
rommem[58] = 33'h101158201;
rommem[59] = 33'h105013382;
rommem[60] = 33'h12AA54830;
rommem[61] = 33'h19768A80A;
rommem[62] = 33'h01A36A5F4;
rommem[63] = 33'h115D034C5;
rommem[64] = 33'h038A53664;
rommem[65] = 33'h1F030C51A;
rommem[66] = 33'h082388505;
rommem[67] = 33'h0203A0148;
rommem[68] = 33'h15082F256;
rommem[69] = 33'h082368501;
rommem[70] = 33'h03664013C;
rommem[71] = 33'h0A5013782;
rommem[72] = 33'h030C51A38;
rommem[73] = 33'h1013DFF10;
rommem[74] = 33'h129823885;
rommem[75] = 33'h0E028A601;
rommem[76] = 33'h142D0FFFF;
rommem[77] = 33'h0D00054C9;
rommem[78] = 33'h00A2AA51A;
rommem[79] = 33'h1E836A6A8;
rommem[80] = 33'h00C1034E4;
rommem[81] = 33'h1050020A9;
rommem[82] = 33'h0E8F49730;
rommem[83] = 33'h1F0D0C8C8;
rommem[84] = 33'h1C9602864;
rommem[85] = 33'h005D00057;
rommem[86] = 33'h0A4822864;
rommem[87] = 33'h00060C900;
rommem[88] = 33'h0FEA906D0;
rommem[89] = 33'h1602885FF;
rommem[90] = 33'h1D00028C9;
rommem[91] = 33'h1FFFDA906;
rommem[92] = 33'h064602885;
rommem[93] = 33'h0FEE06028;
rommem[94] = 33'h16413D0FF;
rommem[95] = 33'h10031C928;
rommem[96] = 33'h1FA8203D0;
rommem[97] = 33'h00030C9FF;
rommem[98] = 33'h1FA8203D0;
rommem[99] = 33'h0FDE060FF;
rommem[100] = 33'h0C90BD0FF;
rommem[101] = 33'h1DBD0001B;
rommem[102] = 33'h185FFFCA9;
rommem[103] = 33'h1FCE06028;
rommem[104] = 33'h0C90BD0FF;
rommem[105] = 33'h0CBD00047;
rommem[106] = 33'h085FFFBA9;
rommem[107] = 33'h0FBE06028;
rommem[108] = 33'h064C0D0FF;
rommem[109] = 33'h10034C928;
rommem[110] = 33'h130A512D0;
rommem[111] = 33'h12A30E2EB;
rommem[112] = 33'h0C22A2A2A;
rommem[113] = 33'h10029EB30;
rommem[114] = 33'h1603085FF;
rommem[115] = 33'h1D00030C9;
rommem[116] = 33'h1BF00A906;
rommem[117] = 33'h1A9603085;
rommem[118] = 33'h03085BF00;
rommem[119] = 33'h0F036A660;
rommem[120] = 33'h00A2AA51F;
rommem[121] = 33'h088F4B7A8;
rommem[122] = 33'h1C8F49788;
rommem[123] = 33'h1E8C8C8C8;
rommem[124] = 33'h1F1D034E4;
rommem[125] = 33'h1050020A9;
rommem[126] = 33'h0C6F49730;
rommem[127] = 33'h000568236;
rommem[128] = 33'h0A536A660;
rommem[129] = 33'h0E8A80A2A;
rommem[130] = 33'h10E1034E4;
rommem[131] = 33'h0B7C8C8CA;
rommem[132] = 33'h0978888F4;
rommem[133] = 33'h1E8C8C8F4;
rommem[134] = 33'h020A9ED80;
rommem[135] = 33'h197300500;
rommem[136] = 33'h136A560F4;
rommem[137] = 33'h1366424F0;
rommem[138] = 33'h036A52C80;
rommem[139] = 33'h11034C51A;
rommem[140] = 33'h08036851D;
rommem[141] = 33'h0F036A521;
rommem[142] = 33'h0F5803A15;
rommem[143] = 33'h00EF038A5;
rommem[144] = 33'h0A507803A;
rommem[145] = 33'h030C51A38;
rommem[146] = 33'h038850410;
rommem[147] = 33'h0A9600880;
rommem[148] = 33'h136640000;
rommem[149] = 33'h0A5483864;
rommem[150] = 33'h1BDAA0A38;
rommem[151] = 33'h06518FA60;
rommem[152] = 33'h1682A8536;
rommem[153] = 33'h00000A060;
rommem[154] = 33'h05A0658A2;
rommem[155] = 33'h034651898;
rommem[156] = 33'h0A8346518;
rommem[157] = 33'h1977AF4B7;
rommem[158] = 33'h1CAC8C8F4;
rommem[159] = 33'h130A5EDD0;
rommem[160] = 33'h0B9A80A3A;
rommem[161] = 33'h1A80AFA60;
rommem[162] = 33'h130A534A6;
rommem[163] = 33'h097002009;
rommem[164] = 33'h1CAC8C8F4;
rommem[165] = 33'h1A960F9D0;
rommem[166] = 33'h0A020000D;
rommem[167] = 33'h1000AA9F2;
rommem[168] = 33'h1DA684858;
rommem[169] = 33'h10000A25A;
rommem[170] = 33'h17A0300FC;
rommem[171] = 33'h13C8560FA;
rommem[172] = 33'h1E2083E86;
rommem[173] = 33'h10000A020;
rommem[174] = 33'h006F03CB7;
rommem[175] = 33'h1C8F2A020;
rommem[176] = 33'h16028F680;
rommem[177] = 33'h0AD5ADA48;
rommem[178] = 33'h1B06AE010;
rommem[179] = 33'h029806A03;
rommem[180] = 33'h0953B40A6;
rommem[181] = 33'h0F2D1A902;
rommem[182] = 33'h002AD0095;
rommem[183] = 33'h0ADFAF0E0;
rommem[184] = 33'h1BDAAE000;
rommem[185] = 33'h0F189F2DF;
rommem[186] = 33'h08DEFF0F2;
rommem[187] = 33'h14085E000;
rommem[188] = 33'h0F2ECA9AA;
rommem[189] = 33'h002B50095;
rommem[190] = 33'h068FA7A1B;
rommem[191] = 33'h18040A540;
rommem[192] = 33'h05ADA48EF;
rommem[193] = 33'h1AA000629;
rommem[194] = 33'h113F30B7C;
rommem[195] = 33'h1F9F35EF3;
rommem[196] = 33'h1DAF2F9F2;
rommem[197] = 33'h10000A25A;
rommem[198] = 33'h0906A44A5;
rommem[199] = 33'h110E0E808;
rommem[200] = 33'h180F7D000;
rommem[201] = 33'h1F38FBDD4;
rommem[202] = 33'h144854405;
rommem[203] = 33'h00029EB8A;
rommem[204] = 33'h0C000090F;
rommem[205] = 33'h0F66918AA;
rommem[206] = 33'h174029500;
rommem[207] = 33'h174FC74FE;
rommem[208] = 33'h0F79568FA;
rommem[209] = 33'h108F89568;
rommem[210] = 33'h08AF69568;
rommem[211] = 33'h10000A968;
rommem[212] = 33'h1A9AA4840;
rommem[213] = 33'h1DF9DF2E1;
rommem[214] = 33'h0008D68F2;
rommem[215] = 33'h0F08A60E0;
rommem[216] = 33'h10840C526;
rommem[217] = 33'h1AAFF0029;
rommem[218] = 33'h195F362A9;
rommem[219] = 33'h1E9388A00;
rommem[220] = 33'h129EBC000;
rommem[221] = 33'h0BDAA000F;
rommem[222] = 33'h0FF49F38F;
rommem[223] = 33'h0854425FF;
rommem[224] = 33'h103D02844;
rommem[225] = 33'h0A9FF5382;
rommem[226] = 33'h004830000;
rommem[227] = 33'h101FF6A82;
rommem[228] = 33'h004000200;
rommem[229] = 33'h010000800;
rommem[230] = 33'h040002000;
rommem[231] = 33'h100008000;
rommem[232] = 33'h000020001;
rommem[233] = 33'h000080004;
rommem[234] = 33'h000200010;
rommem[235] = 33'h0FF800040;
rommem[236] = 33'h0FFFFFFFF;
rommem[237] = 33'h0FFFFFFFF;
rommem[238] = 33'h0FFFFFFFF;
rommem[239] = 33'h0FFFFFFFF;
rommem[240] = 33'h0FFFFFFFF;
rommem[241] = 33'h0FFFFFFFF;
rommem[242] = 33'h0FFFFFFFF;
rommem[243] = 33'h0FFFFFFFF;
rommem[244] = 33'h0FFFFFFFF;
rommem[245] = 33'h0FFFFFFFF;
rommem[246] = 33'h0FFFFFFFF;
rommem[247] = 33'h0FFFFFFFF;
rommem[248] = 33'h0FFFFFFFF;
rommem[249] = 33'h0FFFFFFFF;
rommem[250] = 33'h0FFFFFFFF;
rommem[251] = 33'h0FFFFFFFF;
rommem[252] = 33'h0FFFFFFFF;
rommem[253] = 33'h0FFFFFFFF;
rommem[254] = 33'h0FFFFFFFF;
rommem[255] = 33'h0FFFFFFFF;
rommem[256] = 33'h0FFFFFFFF;
rommem[257] = 33'h0FFFFFFFF;
rommem[258] = 33'h0FFFFFFFF;
rommem[259] = 33'h0FFFFFFFF;
rommem[260] = 33'h0FFFFFFFF;
rommem[261] = 33'h0FFFFFFFF;
rommem[262] = 33'h0FFFFFFFF;
rommem[263] = 33'h0FFFFFFFF;
rommem[264] = 33'h0FFFFFFFF;
rommem[265] = 33'h0FFFFFFFF;
rommem[266] = 33'h0FFFFFFFF;
rommem[267] = 33'h0FFFFFFFF;
rommem[268] = 33'h0FFFFFFFF;
rommem[269] = 33'h0FFFFFFFF;
rommem[270] = 33'h0FFFFFFFF;
rommem[271] = 33'h0FFFFFFFF;
rommem[272] = 33'h0FFFFFFFF;
rommem[273] = 33'h0FFFFFFFF;
rommem[274] = 33'h0FFFFFFFF;
rommem[275] = 33'h0FFFFFFFF;
rommem[276] = 33'h0FFFFFFFF;
rommem[277] = 33'h0FFFFFFFF;
rommem[278] = 33'h0FFFFFFFF;
rommem[279] = 33'h0FFFFFFFF;
rommem[280] = 33'h0FFFFFFFF;
rommem[281] = 33'h0FFFFFFFF;
rommem[282] = 33'h0FFFFFFFF;
rommem[283] = 33'h0FFFFFFFF;
rommem[284] = 33'h0FFFFFFFF;
rommem[285] = 33'h0FFFFFFFF;
rommem[286] = 33'h0FFFFFFFF;
rommem[287] = 33'h0FFFFFFFF;
rommem[288] = 33'h0FFFFFFFF;
rommem[289] = 33'h0FFFFFFFF;
rommem[290] = 33'h0FFFFFFFF;
rommem[291] = 33'h0FFFFFFFF;
rommem[292] = 33'h0FFFFFFFF;
rommem[293] = 33'h0FFFFFFFF;
rommem[294] = 33'h0FFFFFFFF;
rommem[295] = 33'h0FFFFFFFF;
rommem[296] = 33'h0FFFFFFFF;
rommem[297] = 33'h0FFFFFFFF;
rommem[298] = 33'h0FFFFFFFF;
rommem[299] = 33'h0FFFFFFFF;
rommem[300] = 33'h0FFFFFFFF;
rommem[301] = 33'h0FFFFFFFF;
rommem[302] = 33'h0FFFFFFFF;
rommem[303] = 33'h0FFFFFFFF;
rommem[304] = 33'h0FFFFFFFF;
rommem[305] = 33'h0FFFFFFFF;
rommem[306] = 33'h0FFFFFFFF;
rommem[307] = 33'h0FFFFFFFF;
rommem[308] = 33'h0FFFFFFFF;
rommem[309] = 33'h0FFFFFFFF;
rommem[310] = 33'h0FFFFFFFF;
rommem[311] = 33'h0FFFFFFFF;
rommem[312] = 33'h0FFFFFFFF;
rommem[313] = 33'h0FFFFFFFF;
rommem[314] = 33'h0FFFFFFFF;
rommem[315] = 33'h0FFFFFFFF;
rommem[316] = 33'h0FFFFFFFF;
rommem[317] = 33'h0FFFFFFFF;
rommem[318] = 33'h0FFFFFFFF;
rommem[319] = 33'h0FFFFFFFF;
rommem[320] = 33'h0FFFFFFFF;
rommem[321] = 33'h0FFFFFFFF;
rommem[322] = 33'h0FFFFFFFF;
rommem[323] = 33'h0FFFFFFFF;
rommem[324] = 33'h0FFFFFFFF;
rommem[325] = 33'h0FFFFFFFF;
rommem[326] = 33'h0FFFFFFFF;
rommem[327] = 33'h0FFFFFFFF;
rommem[328] = 33'h0FFFFFFFF;
rommem[329] = 33'h0FFFFFFFF;
rommem[330] = 33'h0FFFFFFFF;
rommem[331] = 33'h0FFFFFFFF;
rommem[332] = 33'h0FFFFFFFF;
rommem[333] = 33'h0FFFFFFFF;
rommem[334] = 33'h0FFFFFFFF;
rommem[335] = 33'h0FFFFFFFF;
rommem[336] = 33'h0FFFFFFFF;
rommem[337] = 33'h0FFFFFFFF;
rommem[338] = 33'h0FFFFFFFF;
rommem[339] = 33'h0FFFFFFFF;
rommem[340] = 33'h0FFFFFFFF;
rommem[341] = 33'h0FFFFFFFF;
rommem[342] = 33'h0FFFFFFFF;
rommem[343] = 33'h0FFFFFFFF;
rommem[344] = 33'h0FFFFFFFF;
rommem[345] = 33'h0FFFFFFFF;
rommem[346] = 33'h0FFFFFFFF;
rommem[347] = 33'h0FFFFFFFF;
rommem[348] = 33'h0FFFFFFFF;
rommem[349] = 33'h0FFFFFFFF;
rommem[350] = 33'h0FFFFFFFF;
rommem[351] = 33'h0FFFFFFFF;
rommem[352] = 33'h0FFFFFFFF;
rommem[353] = 33'h0FFFFFFFF;
rommem[354] = 33'h0FFFFFFFF;
rommem[355] = 33'h0FFFFFFFF;
rommem[356] = 33'h0FFFFFFFF;
rommem[357] = 33'h0FFFFFFFF;
rommem[358] = 33'h0FFFFFFFF;
rommem[359] = 33'h0FFFFFFFF;
rommem[360] = 33'h0FFFFFFFF;
rommem[361] = 33'h0FFFFFFFF;
rommem[362] = 33'h0FFFFFFFF;
rommem[363] = 33'h0FFFFFFFF;
rommem[364] = 33'h0FFFFFFFF;
rommem[365] = 33'h0FFFFFFFF;
rommem[366] = 33'h0FFFFFFFF;
rommem[367] = 33'h0FFFFFFFF;
rommem[368] = 33'h0FFFFFFFF;
rommem[369] = 33'h0FFFFFFFF;
rommem[370] = 33'h0FFFFFFFF;
rommem[371] = 33'h0FFFFFFFF;
rommem[372] = 33'h0FFFFFFFF;
rommem[373] = 33'h0FFFFFFFF;
rommem[374] = 33'h0FFFFFFFF;
rommem[375] = 33'h0FFFFFFFF;
rommem[376] = 33'h0FFFFFFFF;
rommem[377] = 33'h0FFFFFFFF;
rommem[378] = 33'h0FFFFFFFF;
rommem[379] = 33'h0FFFFFFFF;
rommem[380] = 33'h0FFFFFFFF;
rommem[381] = 33'h0FFFFFFFF;
rommem[382] = 33'h0FFFFFFFF;
rommem[383] = 33'h0FFFFFFFF;
rommem[384] = 33'h0FFFFFFFF;
rommem[385] = 33'h0FFFFFFFF;
rommem[386] = 33'h0FFFFFFFF;
rommem[387] = 33'h0FFFFFFFF;
rommem[388] = 33'h0FFFFFFFF;
rommem[389] = 33'h0FFFFFFFF;
rommem[390] = 33'h0FFFFFFFF;
rommem[391] = 33'h0FFFFFFFF;
rommem[392] = 33'h0FFFFFFFF;
rommem[393] = 33'h0FFFFFFFF;
rommem[394] = 33'h0FFFFFFFF;
rommem[395] = 33'h0FFFFFFFF;
rommem[396] = 33'h0FFFFFFFF;
rommem[397] = 33'h0FFFFFFFF;
rommem[398] = 33'h0FFFFFFFF;
rommem[399] = 33'h0FFFFFFFF;
rommem[400] = 33'h0FFFFFFFF;
rommem[401] = 33'h0FFFFFFFF;
rommem[402] = 33'h0FFFFFFFF;
rommem[403] = 33'h0FFFFFFFF;
rommem[404] = 33'h0FFFFFFFF;
rommem[405] = 33'h0FFFFFFFF;
rommem[406] = 33'h0FFFFFFFF;
rommem[407] = 33'h0FFFFFFFF;
rommem[408] = 33'h0FFFFFFFF;
rommem[409] = 33'h0FFFFFFFF;
rommem[410] = 33'h0FFFFFFFF;
rommem[411] = 33'h0FFFFFFFF;
rommem[412] = 33'h0FFFFFFFF;
rommem[413] = 33'h0FFFFFFFF;
rommem[414] = 33'h0FFFFFFFF;
rommem[415] = 33'h0FFFFFFFF;
rommem[416] = 33'h0FFFFFFFF;
rommem[417] = 33'h0FFFFFFFF;
rommem[418] = 33'h0FFFFFFFF;
rommem[419] = 33'h0FFFFFFFF;
rommem[420] = 33'h0FFFFFFFF;
rommem[421] = 33'h0FFFFFFFF;
rommem[422] = 33'h0FFFFFFFF;
rommem[423] = 33'h0FFFFFFFF;
rommem[424] = 33'h0FFFFFFFF;
rommem[425] = 33'h0FFFFFFFF;
rommem[426] = 33'h0FFFFFFFF;
rommem[427] = 33'h0FFFFFFFF;
rommem[428] = 33'h0FFFFFFFF;
rommem[429] = 33'h0FFFFFFFF;
rommem[430] = 33'h0FFFFFFFF;
rommem[431] = 33'h0FFFFFFFF;
rommem[432] = 33'h0FFFFFFFF;
rommem[433] = 33'h0FFFFFFFF;
rommem[434] = 33'h0FFFFFFFF;
rommem[435] = 33'h0FFFFFFFF;
rommem[436] = 33'h0FFFFFFFF;
rommem[437] = 33'h0FFFFFFFF;
rommem[438] = 33'h0FFFFFFFF;
rommem[439] = 33'h0FFFFFFFF;
rommem[440] = 33'h0FFFFFFFF;
rommem[441] = 33'h0FFFFFFFF;
rommem[442] = 33'h0FFFFFFFF;
rommem[443] = 33'h0FFFFFFFF;
rommem[444] = 33'h0FFFFFFFF;
rommem[445] = 33'h0FFFFFFFF;
rommem[446] = 33'h0FFFFFFFF;
rommem[447] = 33'h0FFFFFFFF;
rommem[448] = 33'h0FFFFFFFF;
rommem[449] = 33'h0FFFFFFFF;
rommem[450] = 33'h0FFFFFFFF;
rommem[451] = 33'h0FFFFFFFF;
rommem[452] = 33'h0FFFFFFFF;
rommem[453] = 33'h0FFFFFFFF;
rommem[454] = 33'h0FFFFFFFF;
rommem[455] = 33'h0FFFFFFFF;
rommem[456] = 33'h0FFFFFFFF;
rommem[457] = 33'h0FFFFFFFF;
rommem[458] = 33'h0FFFFFFFF;
rommem[459] = 33'h0FFFFFFFF;
rommem[460] = 33'h0FFFFFFFF;
rommem[461] = 33'h0FFFFFFFF;
rommem[462] = 33'h0FFFFFFFF;
rommem[463] = 33'h0FFFFFFFF;
rommem[464] = 33'h0FFFFFFFF;
rommem[465] = 33'h0FFFFFFFF;
rommem[466] = 33'h0FFFFFFFF;
rommem[467] = 33'h0FFFFFFFF;
rommem[468] = 33'h0FFFFFFFF;
rommem[469] = 33'h0FFFFFFFF;
rommem[470] = 33'h0FFFFFFFF;
rommem[471] = 33'h0FFFFFFFF;
rommem[472] = 33'h0FFFFFFFF;
rommem[473] = 33'h0FFFFFFFF;
rommem[474] = 33'h0FFFFFFFF;
rommem[475] = 33'h0FFFFFFFF;
rommem[476] = 33'h0FFFFFFFF;
rommem[477] = 33'h0FFFFFFFF;
rommem[478] = 33'h0FFFFFFFF;
rommem[479] = 33'h0FFFFFFFF;
rommem[480] = 33'h0FFFFFFFF;
rommem[481] = 33'h0FFFFFFFF;
rommem[482] = 33'h0FFFFFFFF;
rommem[483] = 33'h0FFFFFFFF;
rommem[484] = 33'h0FFFFFFFF;
rommem[485] = 33'h0FFFFFFFF;
rommem[486] = 33'h0FFFFFFFF;
rommem[487] = 33'h0FFFFFFFF;
rommem[488] = 33'h0FFFFFFFF;
rommem[489] = 33'h0FFFFFFFF;
rommem[490] = 33'h0FFFFFFFF;
rommem[491] = 33'h0FFFFFFFF;
rommem[492] = 33'h0FFFFFFFF;
rommem[493] = 33'h0FFFFFFFF;
rommem[494] = 33'h0FFFFFFFF;
rommem[495] = 33'h0FFFFFFFF;
rommem[496] = 33'h0FFFFFFFF;
rommem[497] = 33'h0FFFFFFFF;
rommem[498] = 33'h0FFFFFFFF;
rommem[499] = 33'h0FFFFFFFF;
rommem[500] = 33'h0FFFFFFFF;
rommem[501] = 33'h0FFFFFFFF;
rommem[502] = 33'h0FFFFFFFF;
rommem[503] = 33'h0FFFFFFFF;
rommem[504] = 33'h0FFFFFFFF;
rommem[505] = 33'h0FFFFFFFF;
rommem[506] = 33'h0FFFFFFFF;
rommem[507] = 33'h0FFFFFFFF;
rommem[508] = 33'h0FFFFFFFF;
rommem[509] = 33'h0FFFFFFFF;
rommem[510] = 33'h0FFFFFFFF;
rommem[511] = 33'h0FFFFFFFF;
rommem[512] = 33'h06430E208;
rommem[513] = 33'h1FA112009;
rommem[514] = 33'h00A0D0A0D;
rommem[515] = 33'h0646E6553;
rommem[516] = 33'h038353620;
rommem[517] = 33'h063203631;
rommem[518] = 33'h02065646F;
rommem[519] = 33'h149206E69;
rommem[520] = 33'h16C65746E;
rommem[521] = 33'h178654820;
rommem[522] = 33'h1726F6620;
rommem[523] = 33'h12074616D;
rommem[524] = 33'h039207461;
rommem[525] = 33'h030363132;
rommem[526] = 33'h12C6E2C30;
rommem[527] = 33'h020312C38;
rommem[528] = 33'h00A0D3E2D;
rommem[529] = 33'h0A90D6400;
rommem[530] = 33'h1640C8504;
rommem[531] = 33'h1F9C4200B;
rommem[532] = 33'h1F9D03AC9;
rommem[533] = 33'h185F9D020;
rommem[534] = 33'h164088503;
rommem[535] = 33'h0F9D02006;
rommem[536] = 33'h165180585;
rommem[537] = 33'h020088508;
rommem[538] = 33'h10485F9D0;
rommem[539] = 33'h085086518;
rommem[540] = 33'h1F9D02008;
rommem[541] = 33'h065180785;
rommem[542] = 33'h1A5088508;
rommem[543] = 33'h1A62CD007;
rommem[544] = 33'h12000A003;
rommem[545] = 33'h10497F9D0;
rommem[546] = 33'h085086518;
rommem[547] = 33'h1D0CAC808;
rommem[548] = 33'h1F9D020F2;
rommem[549] = 33'h0D0086518;
rommem[550] = 33'h12023A908;
rommem[551] = 33'h0AC82FA05;
rommem[552] = 33'h08546A9FF;
rommem[553] = 33'h1FA052009;
rommem[554] = 33'h1C9FFA282;
rommem[555] = 33'h0C93BF001;
rommem[556] = 33'h1C960F004;
rommem[557] = 33'h02079F005;
rommem[558] = 33'h10A0DFA11;
rommem[559] = 33'h06E550A0D;
rommem[560] = 33'h0776F6E6B;
rommem[561] = 33'h06572206E;
rommem[562] = 33'h164726F63;
rommem[563] = 33'h170797420;
rommem[564] = 33'h100242065;
rommem[565] = 33'h0098507A5;
rommem[566] = 33'h0A9F9F220;
rommem[567] = 33'h0FA05200D;
rommem[568] = 33'h105200AA9;
rommem[569] = 33'h0FF6582FA;
rommem[570] = 33'h1D020B780;
rommem[571] = 33'h1086518F9;
rommem[572] = 33'h111206FF0;
rommem[573] = 33'h00D0A0DFA;
rommem[574] = 33'h06461420A;
rommem[575] = 33'h163657220;
rommem[576] = 33'h02064726F;
rommem[577] = 33'h163656863;
rommem[578] = 33'h06D75736B;
rommem[579] = 33'h1000A0D21;
rommem[580] = 33'h020FEED82;
rommem[581] = 33'h16518F9D0;
rommem[582] = 33'h020088508;
rommem[583] = 33'h00685F9D0;
rommem[584] = 33'h085086518;
rommem[585] = 33'h1F9D02008;
rommem[586] = 33'h0D0086518;
rommem[587] = 33'h0FF1D82BB;
rommem[588] = 33'h018F9D020;
rommem[589] = 33'h108850865;
rommem[590] = 33'h185F9D020;
rommem[591] = 33'h00865180D;
rommem[592] = 33'h0D0200885;
rommem[593] = 33'h1180C85F9;
rommem[594] = 33'h108850865;
rommem[595] = 33'h185F9D020;
rommem[596] = 33'h00865180B;
rommem[597] = 33'h0D0200885;
rommem[598] = 33'h1086518F9;
rommem[599] = 33'h1EC82CDD0;
rommem[600] = 33'h1F009A5FE;
rommem[601] = 33'h1FA11201D;
rommem[602] = 33'h00A0D0A0D;
rommem[603] = 33'h16E776F44;
rommem[604] = 33'h064616F6C;
rommem[605] = 33'h169614620;
rommem[606] = 33'h12E64656C;
rommem[607] = 33'h182000A0D;
rommem[608] = 33'h01120FE7E;
rommem[609] = 33'h00D0A0DFA;
rommem[610] = 33'h0776F440A;
rommem[611] = 33'h0616F6C6E;
rommem[612] = 33'h175532064;
rommem[613] = 33'h173656363;
rommem[614] = 33'h06C756673;
rommem[615] = 33'h04A0A0D21;
rommem[616] = 33'h169706D75;
rommem[617] = 33'h17420676E;
rommem[618] = 33'h10024206F;
rommem[619] = 33'h1F2200DA5;
rommem[620] = 33'h1200CA5F9;
rommem[621] = 33'h00BA5F9F2;
rommem[622] = 33'h120F9F220;
rommem[623] = 33'h10A0DFA11;
rommem[624] = 33'h0000BDC00;
rommem[625] = 33'h0A410C208;
rommem[626] = 33'h0C810B718;
rommem[627] = 33'h060281884;
rommem[628] = 33'h120F9C420;
rommem[629] = 33'h00A0AF9E7;
rommem[630] = 33'h1F0290A0A;
rommem[631] = 33'h1C4200A85;
rommem[632] = 33'h1F9E720F9;
rommem[633] = 33'h0C9600A05;
rommem[634] = 33'h0E902903A;
rommem[635] = 33'h0292FE908;
rommem[636] = 33'h14A48600F;
rommem[637] = 33'h0204A4A4A;
rommem[638] = 33'h12968F9FB;
rommem[639] = 33'h0900AC90F;
rommem[640] = 33'h169066902;
rommem[641] = 33'h110C20830;
rommem[642] = 33'h114971AA4;
rommem[643] = 33'h0281A84C8;
rommem[644] = 33'h000856860;
rommem[645] = 33'h1A0028568;
rommem[646] = 33'h0E600B101;
rommem[647] = 33'h1E602D000;
rommem[648] = 33'h1F0000902;
rommem[649] = 33'h1FA052005;
rommem[650] = 33'h000E6ED80;
rommem[651] = 33'h002E602D0;
rommem[652] = 33'h14300006C;
rommem[653] = 33'h041646F6D;
rommem[654] = 33'h179532037;
rommem[655] = 33'h06D657473;
rommem[656] = 33'h061745320;
rommem[657] = 33'h16E697472;
rommem[658] = 33'h0360A0D67;
rommem[659] = 33'h131384335;
rommem[660] = 33'h06F432036;
rommem[661] = 33'h17461706D;
rommem[662] = 33'h1656C6269;
rommem[663] = 33'h1FF000A0D;
rommem[664] = 33'h1FA620000;
rommem[665] = 33'h0EF26F4C4;
rommem[666] = 33'h1E3EAE988;
rommem[667] = 33'h0D8AEDE4C;
rommem[668] = 33'h1CD72D310;
rommem[669] = 33'h0C236C7D4;
rommem[670] = 33'h1B6FABC98;
rommem[671] = 33'h1ABBEB15C;
rommem[672] = 33'h1A082A620;
rommem[673] = 33'h195469AE4;
rommem[674] = 33'h18A0A8FA8;
rommem[675] = 33'h17ECE846C;
rommem[676] = 33'h173927930;
rommem[677] = 33'h168566DF4;
rommem[678] = 33'h15D1A62B8;
rommem[679] = 33'h0FFFF577C;
rommem[680] = 33'h0FFFFFFFF;
rommem[681] = 33'h0FFFFFFFF;
rommem[682] = 33'h0FFFFFFFF;
rommem[683] = 33'h0FFFFFFFF;
rommem[684] = 33'h0FFFFFFFF;
rommem[685] = 33'h0FFFFFFFF;
rommem[686] = 33'h0FFFFFFFF;
rommem[687] = 33'h0FFFFFFFF;
rommem[688] = 33'h0FFFFFFFF;
rommem[689] = 33'h0FFFFFFFF;
rommem[690] = 33'h0FFFFFFFF;
rommem[691] = 33'h0FFFFFFFF;
rommem[692] = 33'h0FFFFFFFF;
rommem[693] = 33'h0FFFFFFFF;
rommem[694] = 33'h0FFFFFFFF;
rommem[695] = 33'h0FFFFFFFF;
rommem[696] = 33'h0FFFFFFFF;
rommem[697] = 33'h0FFFFFFFF;
rommem[698] = 33'h0FFFFFFFF;
rommem[699] = 33'h0FFFFFFFF;
rommem[700] = 33'h0FFFFFFFF;
rommem[701] = 33'h0FFFFFFFF;
rommem[702] = 33'h0FFFFFFFF;
rommem[703] = 33'h0FFFFFFFF;
rommem[704] = 33'h0FFFFFFFF;
rommem[705] = 33'h0FFFFFFFF;
rommem[706] = 33'h0FFFFFFFF;
rommem[707] = 33'h0FFFFFFFF;
rommem[708] = 33'h0FFFFFFFF;
rommem[709] = 33'h0FFFFFFFF;
rommem[710] = 33'h0FFFFFFFF;
rommem[711] = 33'h0FFFFFFFF;
rommem[712] = 33'h0FFFFFFFF;
rommem[713] = 33'h0FFFFFFFF;
rommem[714] = 33'h0FFFFFFFF;
rommem[715] = 33'h0FFFFFFFF;
rommem[716] = 33'h0FFFFFFFF;
rommem[717] = 33'h0FFFFFFFF;
rommem[718] = 33'h0FFFFFFFF;
rommem[719] = 33'h0FFFFFFFF;
rommem[720] = 33'h0FFFFFFFF;
rommem[721] = 33'h0FFFFFFFF;
rommem[722] = 33'h0FFFFFFFF;
rommem[723] = 33'h0FFFFFFFF;
rommem[724] = 33'h0FFFFFFFF;
rommem[725] = 33'h0FFFFFFFF;
rommem[726] = 33'h0FFFFFFFF;
rommem[727] = 33'h0FFFFFFFF;
rommem[728] = 33'h0FFFFFFFF;
rommem[729] = 33'h0FFFFFFFF;
rommem[730] = 33'h0FFFFFFFF;
rommem[731] = 33'h0FFFFFFFF;
rommem[732] = 33'h0FFFFFFFF;
rommem[733] = 33'h0FFFFFFFF;
rommem[734] = 33'h0FFFFFFFF;
rommem[735] = 33'h0FFFFFFFF;
rommem[736] = 33'h0FFFFFFFF;
rommem[737] = 33'h0FFFFFFFF;
rommem[738] = 33'h0FFFFFFFF;
rommem[739] = 33'h0FFFFFFFF;
rommem[740] = 33'h0FFFFFFFF;
rommem[741] = 33'h0FFFFFFFF;
rommem[742] = 33'h0FFFFFFFF;
rommem[743] = 33'h0FFFFFFFF;
rommem[744] = 33'h0FFFFFFFF;
rommem[745] = 33'h0FFFFFFFF;
rommem[746] = 33'h0FFFFFFFF;
rommem[747] = 33'h0FFFFFFFF;
rommem[748] = 33'h0FFFFFFFF;
rommem[749] = 33'h0FFFFFFFF;
rommem[750] = 33'h0FFFFFFFF;
rommem[751] = 33'h0FFFFFFFF;
rommem[752] = 33'h0FFFFFFFF;
rommem[753] = 33'h0FFFFFFFF;
rommem[754] = 33'h0FFFFFFFF;
rommem[755] = 33'h0FFFFFFFF;
rommem[756] = 33'h0FFFFFFFF;
rommem[757] = 33'h0FFFFFFFF;
rommem[758] = 33'h0FFFFFFFF;
rommem[759] = 33'h0FFFFFFFF;
rommem[760] = 33'h0FFFFFFFF;
rommem[761] = 33'h0FFFFFFFF;
rommem[762] = 33'h0FFFFFFFF;
rommem[763] = 33'h0FFFFFFFF;
rommem[764] = 33'h0FFFFFFFF;
rommem[765] = 33'h0FFFFFFFF;
rommem[766] = 33'h0FFFFFFFF;
rommem[767] = 33'h0FFFFFFFF;
rommem[768] = 33'h0FFFFFFFF;
rommem[769] = 33'h0FFFFFFFF;
rommem[770] = 33'h0FFFFFFFF;
rommem[771] = 33'h0FFFFFFFF;
rommem[772] = 33'h0FFFFFFFF;
rommem[773] = 33'h0FFFFFFFF;
rommem[774] = 33'h0FFFFFFFF;
rommem[775] = 33'h0FFFFFFFF;
rommem[776] = 33'h0FFFFFFFF;
rommem[777] = 33'h0FFFFFFFF;
rommem[778] = 33'h0FFFFFFFF;
rommem[779] = 33'h0FFFFFFFF;
rommem[780] = 33'h0FFFFFFFF;
rommem[781] = 33'h0FFFFFFFF;
rommem[782] = 33'h0FFFFFFFF;
rommem[783] = 33'h0FFFFFFFF;
rommem[784] = 33'h0FFFFFFFF;
rommem[785] = 33'h0FFFFFFFF;
rommem[786] = 33'h0FFFFFFFF;
rommem[787] = 33'h0FFFFFFFF;
rommem[788] = 33'h0FFFFFFFF;
rommem[789] = 33'h0FFFFFFFF;
rommem[790] = 33'h0FFFFFFFF;
rommem[791] = 33'h0FFFFFFFF;
rommem[792] = 33'h0FFFFFFFF;
rommem[793] = 33'h0FFFFFFFF;
rommem[794] = 33'h0FFFFFFFF;
rommem[795] = 33'h0FFFFFFFF;
rommem[796] = 33'h0FFFFFFFF;
rommem[797] = 33'h0FFFFFFFF;
rommem[798] = 33'h0FFFFFFFF;
rommem[799] = 33'h0FFFFFFFF;
rommem[800] = 33'h0FFFFFFFF;
rommem[801] = 33'h0FFFFFFFF;
rommem[802] = 33'h0FFFFFFFF;
rommem[803] = 33'h0FFFFFFFF;
rommem[804] = 33'h0FFFFFFFF;
rommem[805] = 33'h0FFFFFFFF;
rommem[806] = 33'h0FFFFFFFF;
rommem[807] = 33'h0FFFFFFFF;
rommem[808] = 33'h0FFFFFFFF;
rommem[809] = 33'h0FFFFFFFF;
rommem[810] = 33'h0FFFFFFFF;
rommem[811] = 33'h0FFFFFFFF;
rommem[812] = 33'h0FFFFFFFF;
rommem[813] = 33'h0FFFFFFFF;
rommem[814] = 33'h0FFFFFFFF;
rommem[815] = 33'h0FFFFFFFF;
rommem[816] = 33'h0FFFFFFFF;
rommem[817] = 33'h0FFFFFFFF;
rommem[818] = 33'h0FFFFFFFF;
rommem[819] = 33'h0FFFFFFFF;
rommem[820] = 33'h0FFFFFFFF;
rommem[821] = 33'h0FFFFFFFF;
rommem[822] = 33'h0FFFFFFFF;
rommem[823] = 33'h0FFFFFFFF;
rommem[824] = 33'h0FFFFFFFF;
rommem[825] = 33'h0FFFFFFFF;
rommem[826] = 33'h0FFFFFFFF;
rommem[827] = 33'h0FFFFFFFF;
rommem[828] = 33'h0FFFFFFFF;
rommem[829] = 33'h0FFFFFFFF;
rommem[830] = 33'h0FFFFFFFF;
rommem[831] = 33'h0FFFFFFFF;
rommem[832] = 33'h0FFFFFFFF;
rommem[833] = 33'h0FFFFFFFF;
rommem[834] = 33'h0FFFFFFFF;
rommem[835] = 33'h0FFFFFFFF;
rommem[836] = 33'h0FFFFFFFF;
rommem[837] = 33'h0FFFFFFFF;
rommem[838] = 33'h0FFFFFFFF;
rommem[839] = 33'h0FFFFFFFF;
rommem[840] = 33'h0FFFFFFFF;
rommem[841] = 33'h0FFFFFFFF;
rommem[842] = 33'h0FFFFFFFF;
rommem[843] = 33'h0FFFFFFFF;
rommem[844] = 33'h0FFFFFFFF;
rommem[845] = 33'h0FFFFFFFF;
rommem[846] = 33'h0FFFFFFFF;
rommem[847] = 33'h0FFFFFFFF;
rommem[848] = 33'h0FFFFFFFF;
rommem[849] = 33'h0FFFFFFFF;
rommem[850] = 33'h0FFFFFFFF;
rommem[851] = 33'h0FFFFFFFF;
rommem[852] = 33'h0FFFFFFFF;
rommem[853] = 33'h0FFFFFFFF;
rommem[854] = 33'h0FFFFFFFF;
rommem[855] = 33'h0FFFFFFFF;
rommem[856] = 33'h0FFFFFFFF;
rommem[857] = 33'h0FFFFFFFF;
rommem[858] = 33'h0FFFFFFFF;
rommem[859] = 33'h0FFFFFFFF;
rommem[860] = 33'h0FFFFFFFF;
rommem[861] = 33'h0FFFFFFFF;
rommem[862] = 33'h0FFFFFFFF;
rommem[863] = 33'h0FFFFFFFF;
rommem[864] = 33'h0FFFFFFFF;
rommem[865] = 33'h0FFFFFFFF;
rommem[866] = 33'h0FFFFFFFF;
rommem[867] = 33'h0FFFFFFFF;
rommem[868] = 33'h0FFFFFFFF;
rommem[869] = 33'h0FFFFFFFF;
rommem[870] = 33'h0FFFFFFFF;
rommem[871] = 33'h0FFFFFFFF;
rommem[872] = 33'h0FFFFFFFF;
rommem[873] = 33'h0FFFFFFFF;
rommem[874] = 33'h0FFFFFFFF;
rommem[875] = 33'h0FFFFFFFF;
rommem[876] = 33'h0FFFFFFFF;
rommem[877] = 33'h0FFFFFFFF;
rommem[878] = 33'h0FFFFFFFF;
rommem[879] = 33'h0FFFFFFFF;
rommem[880] = 33'h0FFFFFFFF;
rommem[881] = 33'h0FFFFFFFF;
rommem[882] = 33'h0FFFFFFFF;
rommem[883] = 33'h0FFFFFFFF;
rommem[884] = 33'h0FFFFFFFF;
rommem[885] = 33'h0FFFFFFFF;
rommem[886] = 33'h0FFFFFFFF;
rommem[887] = 33'h0FFFFFFFF;
rommem[888] = 33'h0FFFFFFFF;
rommem[889] = 33'h0FFFFFFFF;
rommem[890] = 33'h0FFFFFFFF;
rommem[891] = 33'h0FFFFFFFF;
rommem[892] = 33'h0FFFFFFFF;
rommem[893] = 33'h0FFFFFFFF;
rommem[894] = 33'h0FFFFFFFF;
rommem[895] = 33'h0FFFFFFFF;
rommem[896] = 33'h0FFFFFFFF;
rommem[897] = 33'h0FFFFFFFF;
rommem[898] = 33'h0FFFFFFFF;
rommem[899] = 33'h0FFFFFFFF;
rommem[900] = 33'h0FFFFFFFF;
rommem[901] = 33'h0FFFFFFFF;
rommem[902] = 33'h0FFFFFFFF;
rommem[903] = 33'h0FFFFFFFF;
rommem[904] = 33'h0FFFFFFFF;
rommem[905] = 33'h0FFFFFFFF;
rommem[906] = 33'h0FFFFFFFF;
rommem[907] = 33'h0FFFFFFFF;
rommem[908] = 33'h0FFFFFFFF;
rommem[909] = 33'h0FFFFFFFF;
rommem[910] = 33'h0FFFFFFFF;
rommem[911] = 33'h0FFFFFFFF;
rommem[912] = 33'h0FFFFFFFF;
rommem[913] = 33'h0FFFFFFFF;
rommem[914] = 33'h0FFFFFFFF;
rommem[915] = 33'h0FFFFFFFF;
rommem[916] = 33'h0FFFFFFFF;
rommem[917] = 33'h0FFFFFFFF;
rommem[918] = 33'h0FFFFFFFF;
rommem[919] = 33'h0FFFFFFFF;
rommem[920] = 33'h0FFFFFFFF;
rommem[921] = 33'h0FFFFFFFF;
rommem[922] = 33'h0FFFFFFFF;
rommem[923] = 33'h0FFFFFFFF;
rommem[924] = 33'h0FFFFFFFF;
rommem[925] = 33'h0FFFFFFFF;
rommem[926] = 33'h0FFFFFFFF;
rommem[927] = 33'h0FFFFFFFF;
rommem[928] = 33'h0FFFFFFFF;
rommem[929] = 33'h0FFFFFFFF;
rommem[930] = 33'h0FFFFFFFF;
rommem[931] = 33'h0FFFFFFFF;
rommem[932] = 33'h0FFFFFFFF;
rommem[933] = 33'h0FFFFFFFF;
rommem[934] = 33'h0FFFFFFFF;
rommem[935] = 33'h0FFFFFFFF;
rommem[936] = 33'h0FFFFFFFF;
rommem[937] = 33'h0FFFFFFFF;
rommem[938] = 33'h0FFFFFFFF;
rommem[939] = 33'h0FFFFFFFF;
rommem[940] = 33'h0FFFFFFFF;
rommem[941] = 33'h0FFFFFFFF;
rommem[942] = 33'h0FFFFFFFF;
rommem[943] = 33'h0FFFFFFFF;
rommem[944] = 33'h0FFFFFFFF;
rommem[945] = 33'h0FFFFFFFF;
rommem[946] = 33'h0FFFFFFFF;
rommem[947] = 33'h0FFFFFFFF;
rommem[948] = 33'h0FFFFFFFF;
rommem[949] = 33'h0FFFFFFFF;
rommem[950] = 33'h0FFFFFFFF;
rommem[951] = 33'h0FFFFFFFF;
rommem[952] = 33'h0FFFFFFFF;
rommem[953] = 33'h0FFFFFFFF;
rommem[954] = 33'h0FFFFFFFF;
rommem[955] = 33'h0FFFFFFFF;
rommem[956] = 33'h0FFFFFFFF;
rommem[957] = 33'h0FFFFFFFF;
rommem[958] = 33'h0FFFFFFFF;
rommem[959] = 33'h0FFFFFFFF;
rommem[960] = 33'h0FFFFFFFF;
rommem[961] = 33'h0FFFFFFFF;
rommem[962] = 33'h0FFFFFFFF;
rommem[963] = 33'h0FFFFFFFF;
rommem[964] = 33'h0FFFFFFFF;
rommem[965] = 33'h0FFFFFFFF;
rommem[966] = 33'h0FFFFFFFF;
rommem[967] = 33'h0FFFFFFFF;
rommem[968] = 33'h0FFFFFFFF;
rommem[969] = 33'h0FFFFFFFF;
rommem[970] = 33'h0FFFFFFFF;
rommem[971] = 33'h0FFFFFFFF;
rommem[972] = 33'h0FFFFFFFF;
rommem[973] = 33'h0FFFFFFFF;
rommem[974] = 33'h0FFFFFFFF;
rommem[975] = 33'h0FFFFFFFF;
rommem[976] = 33'h0FFFFFFFF;
rommem[977] = 33'h0FFFFFFFF;
rommem[978] = 33'h0FFFFFFFF;
rommem[979] = 33'h0FFFFFFFF;
rommem[980] = 33'h0FFFFFFFF;
rommem[981] = 33'h0FFFFFFFF;
rommem[982] = 33'h0FFFFFFFF;
rommem[983] = 33'h0FFFFFFFF;
rommem[984] = 33'h0FFFFFFFF;
rommem[985] = 33'h0FFFFFFFF;
rommem[986] = 33'h0FFFFFFFF;
rommem[987] = 33'h0FFFFFFFF;
rommem[988] = 33'h0FFFFFFFF;
rommem[989] = 33'h0FFFFFFFF;
rommem[990] = 33'h0FFFFFFFF;
rommem[991] = 33'h0FFFFFFFF;
rommem[992] = 33'h0FFFFFFFF;
rommem[993] = 33'h0FFFFFFFF;
rommem[994] = 33'h0FFFFFFFF;
rommem[995] = 33'h0FFFFFFFF;
rommem[996] = 33'h0FFFFFFFF;
rommem[997] = 33'h0FFFFFFFF;
rommem[998] = 33'h0FFFFFFFF;
rommem[999] = 33'h0FFFFFFFF;
rommem[1000] = 33'h0FFFFFFFF;
rommem[1001] = 33'h0FFFFFFFF;
rommem[1002] = 33'h0FFFFFFFF;
rommem[1003] = 33'h0FFFFFFFF;
rommem[1004] = 33'h0FFFFFFFF;
rommem[1005] = 33'h0FFFFFFFF;
rommem[1006] = 33'h0FFFFFFFF;
rommem[1007] = 33'h0FFFFFFFF;
rommem[1008] = 33'h0FFFFFFFF;
rommem[1009] = 33'h0FFFFFFFF;
rommem[1010] = 33'h0FFFFFFFF;
rommem[1011] = 33'h0FFFFFFFF;
rommem[1012] = 33'h0FFFFFFFF;
rommem[1013] = 33'h0FFFFFFFF;
rommem[1014] = 33'h0FFFFFFFF;
rommem[1015] = 33'h0FFFFFFFF;
rommem[1016] = 33'h0FFFFFFFF;
rommem[1017] = 33'h0FFFFFFFF;
rommem[1018] = 33'h0FFFFFFFF;
rommem[1019] = 33'h0FFFFFFFF;
rommem[1020] = 33'h0FFFFFFFF;
rommem[1021] = 33'h0FFFFFFFF;
rommem[1022] = 33'h0FFFFFFFF;
rommem[1023] = 33'h0F06CF000;
