/*
ORSoC GFX accelerator core
Copyright 2012, ORSoC, Per Lenander, Anton Fosselius.

PER-PIXEL COLORING MODULE

 This file is part of orgfx.

 orgfx is free software: you can redistribute it and/or modify
 it under the terms of the GNU Lesser General Public License as published by
 the Free Software Foundation, either version 3 of the License, or
 (at your option) any later version. 

 orgfx is distributed in the hope that it will be useful,
 but WITHOUT ANY WARRANTY; without even the implied warranty of
 MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 GNU Lesser General Public License for more details.

 You should have received a copy of the GNU Lesser General Public License
 along with orgfx.  If not, see <http://www.gnu.org/licenses/>.

 Robert Finch
 Modified to support greater number of color depths.
*/

/*
This module adds color to the pixel generated by the rasterizer. It can either draw a flat color (using pixel_color_i) or
colors from a texture by using the u and v coordinates generated by the rasterizer. 
*/
module gfx_fragment_processor(clk_i, rst_i,
  pixel_alpha_i,
  x_counter_i, y_counter_i, z_i, u_i, v_i, bezier_factor0_i, bezier_factor1_i, bezier_inside_i, write_i, curve_write_i, ack_o, // from raster
  pixel_x_o, pixel_y_o, pixel_z_o, pixel_color_i, pixel_color_o, pixel_alpha_o, write_o, ack_i,  // to blender
  texture_ack_i, texture_data_i, texture_addr_o, texture_request_o, // to/from wishbone master read
  texture_enable_i, tex0_base_i, tex0_size_x_i, tex0_size_y_i, color_depth_i, colorkey_enable_i, colorkey_i // from wishbone slave
  );

parameter point_width = 16;

input clk_i;
input rst_i;

input [7:0]  pixel_alpha_i;

// from raster
input [point_width-1:0] x_counter_i;
input [point_width-1:0] y_counter_i;
input signed [point_width-1:0] z_i;
input [point_width-1:0] u_i; // x-ish texture coordinate
input [point_width-1:0] v_i; // y-ish texture coordinate
input [point_width-1:0] bezier_factor0_i; // Used for curve writing
input [point_width-1:0] bezier_factor1_i; // Used for curve writing
input                   bezier_inside_i;
input            [31:0] pixel_color_i;
input                   write_i;
input                   curve_write_i;
output reg              ack_o;

//to render
output reg [point_width-1:0] pixel_x_o;
output reg [point_width-1:0] pixel_y_o;
output reg signed [point_width-1:0] pixel_z_o;
output reg            [31:0] pixel_color_o;
output reg             [7:0] pixel_alpha_o;
output reg                   write_o;
input                        ack_i;

// to/from wishbone master read
input              texture_ack_i;
input      [127:0] texture_data_i;
output      [31:0] texture_addr_o;
output reg         texture_request_o;

// from wishbone slave
input                   texture_enable_i;
input            [31:2] tex0_base_i;
input [point_width-1:0] tex0_size_x_i;
input [point_width-1:0] tex0_size_y_i;
input            [ 1:0] color_depth_i;
input                   colorkey_enable_i;
input            [31:0] colorkey_i;

wire             [31:0] pixel_offset;

// Calculate the memory address of the texel to read 
wire [6:0] mb, me;

gfx_CalcAddress u1
(
	.base_address_i(tex0_base_i),
	.color_depth_i(color_depth_i),
	.hdisplayed_i(tex0_size_x_i),
	.x_coord_i(u_i),
	.y_coord_i(v_i),
	.address_o(texture_addr_o),
	.mb_o(mb),
	.me_o(me)
);

// State machine
reg [1:0] state;
parameter wait_state = 2'b00, texture_read_state = 2'b01, write_pixel_state = 2'b10;

parameter BPP6 = 3'd0;
parameter BPP8 = 3'd1;
parameter BPP9 = 3'd2;
parameter BPP12 = 3'd3;
parameter BPP15 = 3'd4;
parameter BPP16 = 3'd5;
parameter BPP24 = 3'd6;
parameter BPP32 = 3'd7;

wire [31:0] mem_conv_color_o;

// Color converter
memory_to_color memory_proc(
.mem_i (texture_data_i),
.mb_i (mb),
.me_i (me),
.color_o (mem_conv_color_o)
);

// Does the fetched texel match the colorkey?
reg transparent_pixel;
always @(color_depth_i or mem_conv_color_o or colorkey_i)
case(color_depth_i)
BPP6:	transparent_pixel = mem_conv_color_o[5:0] == colorkey_i[5:0];
BPP8:	transparent_pixel = mem_conv_color_o[7:0] == colorkey_i[7:0];
BPP9:	transparent_pixel = mem_conv_color_o[8:0] == colorkey_i[8:0];
BPP12:	transparent_pixel = mem_conv_color_o[11:0] == colorkey_i[11:0];
BPP15:	transparent_pixel = mem_conv_color_o[14:0] == colorkey_i[14:0];
BPP16:	transparent_pixel = mem_conv_color_o[15:0] == colorkey_i[15:0];
BPP24:	transparent_pixel = mem_conv_color_o[23:0] == colorkey_i[23:0];
BPP32:	transparent_pixel = mem_conv_color_o[23:0] == colorkey_i[23:0];
endcase

// These variables are used when rendering bezier shapes. If bezier_draw is true, pixel is drawn, if it is false, pixel is discarded.
// These variables are only used if curve_write_i is high

// Calculate if factor0*factor0 > factor1
// Values are in the range [0..1], represented by a [point_width-1:0] bit array
wire [2*point_width-1:0] bezier_factor0_squared = bezier_factor0_i*bezier_factor0_i;
wire bezier_eval = bezier_factor0_squared[2*point_width-1:point_width] > bezier_factor1_i;
wire bezier_draw = bezier_inside_i ^ bezier_eval; // inside xor eval

// Acknowledge when a command has completed
always @(posedge clk_i or posedge rst_i)
begin
  // reset, init component
  if(rst_i)
  begin
    ack_o             <= 1'b0;
    write_o           <= 1'b0;
    pixel_x_o         <= 1'b0;
    pixel_y_o         <= 1'b0;
    pixel_z_o         <= 1'b0;
    pixel_color_o     <= 1'b0;
    pixel_alpha_o     <= 1'b0;
    texture_request_o <= 1'b0;
  end
  // Else, set outputs for next cycle
  else
  begin
    case (state)

      wait_state:
      begin
        ack_o   <= write_i & curve_write_i & ~bezier_draw;

        if(write_i & texture_enable_i & (~curve_write_i | bezier_draw))
          texture_request_o <= 1'b1;
        else if(write_i & (~curve_write_i | bezier_draw))
        begin
          pixel_x_o         <= x_counter_i;
          pixel_y_o         <= y_counter_i;
          pixel_z_o         <= z_i;
          pixel_color_o     <= pixel_color_i;
          pixel_alpha_o     <= pixel_alpha_i;
          write_o           <= 1'b1; // Note, colorkey only supported for texture reads
        end
      end


      texture_read_state:
        if(texture_ack_i)
        begin
          pixel_x_o         <= x_counter_i;
          pixel_y_o         <= y_counter_i;
          pixel_z_o         <= z_i;
          pixel_color_o     <= mem_conv_color_o;
          pixel_alpha_o     <= pixel_alpha_i;
          texture_request_o <= 1'b0;
          if(colorkey_enable_i & transparent_pixel)
            ack_o           <= 1'b1; // Colorkey enabled: Only write if the pixel doesn't match the colorkey
          else
            write_o         <= 1'b1;
        end


      write_pixel_state:
      begin
        write_o  <= 1'b0;
        ack_o    <= ack_i;
      end

    endcase
  end
end

// State machine
always @(posedge clk_i or posedge rst_i)
begin
  // reset, init component
  if(rst_i)
    state <= wait_state;
  // Move in statemachine
  else
    case (state)

      wait_state:
        if(write_i & texture_enable_i & (~curve_write_i | bezier_draw))
          state <= texture_read_state;
        else if(write_i & (~curve_write_i | bezier_draw))
          state <= write_pixel_state;

      texture_read_state:
        // Check for texture ack. If we have colorkeying enabled, only goto the write state if the texture doesn't match the colorkey
        if(texture_ack_i & colorkey_enable_i)
          state <= transparent_pixel ? wait_state : write_pixel_state;
        else if(texture_ack_i)
          state <= write_pixel_state;

      write_pixel_state:
        if(ack_i)
          state <= wait_state;

    endcase
end

endmodule

