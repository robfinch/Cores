XCHG_MEM:
begin
	res <= b;
	tGoto(STORE_DATA);
end
