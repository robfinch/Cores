RsqrteLUT[0] = 32'h3f800000;
RsqrteLUT[1] = 32'h42000000;
RsqrteLUT[2] = 32'h41b504f3;
RsqrteLUT[3] = 32'h4193cd3a;
RsqrteLUT[4] = 32'h41800000;
RsqrteLUT[5] = 32'h4164f92e;
RsqrteLUT[6] = 32'h415105eb;
RsqrteLUT[7] = 32'h4141848f;
RsqrteLUT[8] = 32'h413504f3;
RsqrteLUT[9] = 32'h412aaaaa;
RsqrteLUT[10] = 32'h4121e89b;
RsqrteLUT[11] = 32'h411a5fb1;
RsqrteLUT[12] = 32'h4113cd3a;
RsqrteLUT[13] = 32'h410e00d5;
RsqrteLUT[14] = 32'h4108d677;
RsqrteLUT[15] = 32'h410432a5;
RsqrteLUT[16] = 32'h41000000;
RsqrteLUT[17] = 32'h40f85b42;
RsqrteLUT[18] = 32'h40f15bee;
RsqrteLUT[19] = 32'h40eaebf5;
RsqrteLUT[20] = 32'h40e4f92e;
RsqrteLUT[21] = 32'h40df7482;
RsqrteLUT[22] = 32'h40da5149;
RsqrteLUT[23] = 32'h40d584cd;
RsqrteLUT[24] = 32'h40d105eb;
RsqrteLUT[25] = 32'h40cccccc;
RsqrteLUT[26] = 32'h40c8d2ab;
RsqrteLUT[27] = 32'h40c511a2;
RsqrteLUT[28] = 32'h40c1848f;
RsqrteLUT[29] = 32'h40be26eb;
RsqrteLUT[30] = 32'h40baf4ba;
RsqrteLUT[31] = 32'h40b7ea73;
RsqrteLUT[32] = 32'h40b504f3;
RsqrteLUT[33] = 32'h40b24169;
RsqrteLUT[34] = 32'h40af9d53;
RsqrteLUT[35] = 32'h40ad166c;
RsqrteLUT[36] = 32'h40aaaaaa;
RsqrteLUT[37] = 32'h40a85835;
RsqrteLUT[38] = 32'h40a61d5f;
RsqrteLUT[39] = 32'h40a3f8a2;
RsqrteLUT[40] = 32'h40a1e89b;
RsqrteLUT[41] = 32'h409fec03;
RsqrteLUT[42] = 32'h409e01b2;
RsqrteLUT[43] = 32'h409c2895;
RsqrteLUT[44] = 32'h409a5fb1;
RsqrteLUT[45] = 32'h4098a61e;
RsqrteLUT[46] = 32'h4096fb06;
RsqrteLUT[47] = 32'h40955da1;
RsqrteLUT[48] = 32'h4093cd3a;
RsqrteLUT[49] = 32'h40924924;
RsqrteLUT[50] = 32'h4090d0c2;
RsqrteLUT[51] = 32'h408f6380;
RsqrteLUT[52] = 32'h408e00d5;
RsqrteLUT[53] = 32'h408ca83f;
RsqrteLUT[54] = 32'h408b5947;
RsqrteLUT[55] = 32'h408a137d;
RsqrteLUT[56] = 32'h4088d677;
RsqrteLUT[57] = 32'h4087a1d2;
RsqrteLUT[58] = 32'h40867531;
RsqrteLUT[59] = 32'h4085503d;
RsqrteLUT[60] = 32'h408432a5;
RsqrteLUT[61] = 32'h40831c19;
RsqrteLUT[62] = 32'h40820c52;
RsqrteLUT[63] = 32'h4081030a;
RsqrteLUT[64] = 32'h40800000;
RsqrteLUT[65] = 32'h407e05ec;
RsqrteLUT[66] = 32'h407c1764;
RsqrteLUT[67] = 32'h407a33f9;
RsqrteLUT[68] = 32'h40785b42;
RsqrteLUT[69] = 32'h40768cdb;
RsqrteLUT[70] = 32'h4074c866;
RsqrteLUT[71] = 32'h40730d89;
RsqrteLUT[72] = 32'h40715bee;
RsqrteLUT[73] = 32'h406fb344;
RsqrteLUT[74] = 32'h406e133d;
RsqrteLUT[75] = 32'h406c7b90;
RsqrteLUT[76] = 32'h406aebf5;
RsqrteLUT[77] = 32'h40696429;
RsqrteLUT[78] = 32'h4067e3ed;
RsqrteLUT[79] = 32'h40666b02;
RsqrteLUT[80] = 32'h4064f92e;
RsqrteLUT[81] = 32'h40638e38;
RsqrteLUT[82] = 32'h406229ec;
RsqrteLUT[83] = 32'h4060cc15;
RsqrteLUT[84] = 32'h405f7482;
RsqrteLUT[85] = 32'h405e2304;
RsqrteLUT[86] = 32'h405cd76d;
RsqrteLUT[87] = 32'h405b9192;
RsqrteLUT[88] = 32'h405a5149;
RsqrteLUT[89] = 32'h4059166a;
RsqrteLUT[90] = 32'h4057e0ce;
RsqrteLUT[91] = 32'h4056b050;
RsqrteLUT[92] = 32'h405584cd;
RsqrteLUT[93] = 32'h40545e22;
RsqrteLUT[94] = 32'h40533c2d;
RsqrteLUT[95] = 32'h40521ed0;
RsqrteLUT[96] = 32'h405105eb;
RsqrteLUT[97] = 32'h404ff161;
RsqrteLUT[98] = 32'h404ee115;
RsqrteLUT[99] = 32'h404dd4ed;
RsqrteLUT[100] = 32'h404ccccc;
RsqrteLUT[101] = 32'h404bc89b;
RsqrteLUT[102] = 32'h404ac83f;
RsqrteLUT[103] = 32'h4049cba1;
RsqrteLUT[104] = 32'h4048d2ab;
RsqrteLUT[105] = 32'h4047dd45;
RsqrteLUT[106] = 32'h4046eb5a;
RsqrteLUT[107] = 32'h4045fcd5;
RsqrteLUT[108] = 32'h404511a2;
RsqrteLUT[109] = 32'h404429ae;
RsqrteLUT[110] = 32'h404344e6;
RsqrteLUT[111] = 32'h40426336;
RsqrteLUT[112] = 32'h4041848f;
RsqrteLUT[113] = 32'h4040a8dd;
RsqrteLUT[114] = 32'h403fd011;
RsqrteLUT[115] = 32'h403efa1b;
RsqrteLUT[116] = 32'h403e26eb;
RsqrteLUT[117] = 32'h403d5671;
RsqrteLUT[118] = 32'h403c889f;
RsqrteLUT[119] = 32'h403bbd66;
RsqrteLUT[120] = 32'h403af4ba;
RsqrteLUT[121] = 32'h403a2e8b;
RsqrteLUT[122] = 32'h40396ace;
RsqrteLUT[123] = 32'h4038a974;
RsqrteLUT[124] = 32'h4037ea73;
RsqrteLUT[125] = 32'h40372dbe;
RsqrteLUT[126] = 32'h40367349;
RsqrteLUT[127] = 32'h4035bb09;
RsqrteLUT[128] = 32'h403504f3;
RsqrteLUT[129] = 32'h403450fc;
RsqrteLUT[130] = 32'h40339f19;
RsqrteLUT[131] = 32'h4032ef41;
RsqrteLUT[132] = 32'h40324169;
RsqrteLUT[133] = 32'h40319589;
RsqrteLUT[134] = 32'h4030eb95;
RsqrteLUT[135] = 32'h40304386;
RsqrteLUT[136] = 32'h402f9d53;
RsqrteLUT[137] = 32'h402ef8f2;
RsqrteLUT[138] = 32'h402e565b;
RsqrteLUT[139] = 32'h402db587;
RsqrteLUT[140] = 32'h402d166c;
RsqrteLUT[141] = 32'h402c7903;
RsqrteLUT[142] = 32'h402bdd45;
RsqrteLUT[143] = 32'h402b432a;
RsqrteLUT[144] = 32'h402aaaaa;
RsqrteLUT[145] = 32'h402a13bf;
RsqrteLUT[146] = 32'h40297e62;
RsqrteLUT[147] = 32'h4028ea8b;
RsqrteLUT[148] = 32'h40285835;
RsqrteLUT[149] = 32'h4027c758;
RsqrteLUT[150] = 32'h402737ef;
RsqrteLUT[151] = 32'h4026a9f3;
RsqrteLUT[152] = 32'h40261d5f;
RsqrteLUT[153] = 32'h4025922c;
RsqrteLUT[154] = 32'h40250854;
RsqrteLUT[155] = 32'h40247fd3;
RsqrteLUT[156] = 32'h4023f8a2;
RsqrteLUT[157] = 32'h402372bc;
RsqrteLUT[158] = 32'h4022ee1d;
RsqrteLUT[159] = 32'h40226abe;
RsqrteLUT[160] = 32'h4021e89b;
RsqrteLUT[161] = 32'h402167ae;
RsqrteLUT[162] = 32'h4020e7f4;
RsqrteLUT[163] = 32'h40206967;
RsqrteLUT[164] = 32'h401fec03;
RsqrteLUT[165] = 32'h401f6fc3;
RsqrteLUT[166] = 32'h401ef4a4;
RsqrteLUT[167] = 32'h401e7a9f;
RsqrteLUT[168] = 32'h401e01b2;
RsqrteLUT[169] = 32'h401d89d8;
RsqrteLUT[170] = 32'h401d130d;
RsqrteLUT[171] = 32'h401c9d4e;
RsqrteLUT[172] = 32'h401c2895;
RsqrteLUT[173] = 32'h401bb4e0;
RsqrteLUT[174] = 32'h401b422b;
RsqrteLUT[175] = 32'h401ad072;
RsqrteLUT[176] = 32'h401a5fb1;
RsqrteLUT[177] = 32'h4019efe6;
RsqrteLUT[178] = 32'h4019810c;
RsqrteLUT[179] = 32'h4019131f;
RsqrteLUT[180] = 32'h4018a61e;
RsqrteLUT[181] = 32'h40183a05;
RsqrteLUT[182] = 32'h4017cecf;
RsqrteLUT[183] = 32'h4017647b;
RsqrteLUT[184] = 32'h4016fb06;
RsqrteLUT[185] = 32'h4016926b;
RsqrteLUT[186] = 32'h40162aa9;
RsqrteLUT[187] = 32'h4015c3bc;
RsqrteLUT[188] = 32'h40155da1;
RsqrteLUT[189] = 32'h4014f857;
RsqrteLUT[190] = 32'h401493d9;
RsqrteLUT[191] = 32'h40143025;
RsqrteLUT[192] = 32'h4013cd3a;
RsqrteLUT[193] = 32'h40136b13;
RsqrteLUT[194] = 32'h401309af;
RsqrteLUT[195] = 32'h4012a90b;
RsqrteLUT[196] = 32'h40124924;
RsqrteLUT[197] = 32'h4011e9f9;
RsqrteLUT[198] = 32'h40118b86;
RsqrteLUT[199] = 32'h40112dca;
RsqrteLUT[200] = 32'h4010d0c2;
RsqrteLUT[201] = 32'h4010746c;
RsqrteLUT[202] = 32'h401018c6;
RsqrteLUT[203] = 32'h400fbdcd;
RsqrteLUT[204] = 32'h400f6380;
RsqrteLUT[205] = 32'h400f09dc;
RsqrteLUT[206] = 32'h400eb0e0;
RsqrteLUT[207] = 32'h400e5888;
RsqrteLUT[208] = 32'h400e00d5;
RsqrteLUT[209] = 32'h400da9c2;
RsqrteLUT[210] = 32'h400d534f;
RsqrteLUT[211] = 32'h400cfd79;
RsqrteLUT[212] = 32'h400ca83f;
RsqrteLUT[213] = 32'h400c539f;
RsqrteLUT[214] = 32'h400bff97;
RsqrteLUT[215] = 32'h400bac25;
RsqrteLUT[216] = 32'h400b5947;
RsqrteLUT[217] = 32'h400b06fd;
RsqrteLUT[218] = 32'h400ab543;
RsqrteLUT[219] = 32'h400a6419;
RsqrteLUT[220] = 32'h400a137d;
RsqrteLUT[221] = 32'h4009c36d;
RsqrteLUT[222] = 32'h400973e8;
RsqrteLUT[223] = 32'h400924eb;
RsqrteLUT[224] = 32'h4008d677;
RsqrteLUT[225] = 32'h40088888;
RsqrteLUT[226] = 32'h40083b1e;
RsqrteLUT[227] = 32'h4007ee37;
RsqrteLUT[228] = 32'h4007a1d2;
RsqrteLUT[229] = 32'h400755ed;
RsqrteLUT[230] = 32'h40070a86;
RsqrteLUT[231] = 32'h4006bf9e;
RsqrteLUT[232] = 32'h40067531;
RsqrteLUT[233] = 32'h40062b3f;
RsqrteLUT[234] = 32'h4005e1c7;
RsqrteLUT[235] = 32'h400598c7;
RsqrteLUT[236] = 32'h4005503d;
RsqrteLUT[237] = 32'h4005082a;
RsqrteLUT[238] = 32'h4004c08b;
RsqrteLUT[239] = 32'h4004795f;
RsqrteLUT[240] = 32'h400432a5;
RsqrteLUT[241] = 32'h4003ec5b;
RsqrteLUT[242] = 32'h4003a682;
RsqrteLUT[243] = 32'h40036117;
RsqrteLUT[244] = 32'h40031c19;
RsqrteLUT[245] = 32'h4002d788;
RsqrteLUT[246] = 32'h40029361;
RsqrteLUT[247] = 32'h40024fa5;
RsqrteLUT[248] = 32'h40020c52;
RsqrteLUT[249] = 32'h4001c966;
RsqrteLUT[250] = 32'h400186e2;
RsqrteLUT[251] = 32'h400144c3;
RsqrteLUT[252] = 32'h4001030a;
RsqrteLUT[253] = 32'h4000c1b4;
RsqrteLUT[254] = 32'h400080c1;
RsqrteLUT[255] = 32'h40004030;
RsqrteLUT[256] = 32'h40000000;
RsqrteLUT[257] = 32'h3fff805f;
RsqrteLUT[258] = 32'h3fff017d;
RsqrteLUT[259] = 32'h3ffe8357;
RsqrteLUT[260] = 32'h3ffe05ec;
RsqrteLUT[261] = 32'h3ffd8939;
RsqrteLUT[262] = 32'h3ffd0d3d;
RsqrteLUT[263] = 32'h3ffc91f7;
RsqrteLUT[264] = 32'h3ffc1764;
RsqrteLUT[265] = 32'h3ffb9d82;
RsqrteLUT[266] = 32'h3ffb2451;
RsqrteLUT[267] = 32'h3ffaabcf;
RsqrteLUT[268] = 32'h3ffa33f9;
RsqrteLUT[269] = 32'h3ff9bcce;
RsqrteLUT[270] = 32'h3ff9464d;
RsqrteLUT[271] = 32'h3ff8d074;
RsqrteLUT[272] = 32'h3ff85b42;
RsqrteLUT[273] = 32'h3ff7e6b4;
RsqrteLUT[274] = 32'h3ff772ca;
RsqrteLUT[275] = 32'h3ff6ff83;
RsqrteLUT[276] = 32'h3ff68cdb;
RsqrteLUT[277] = 32'h3ff61ad3;
RsqrteLUT[278] = 32'h3ff5a968;
RsqrteLUT[279] = 32'h3ff5389a;
RsqrteLUT[280] = 32'h3ff4c866;
RsqrteLUT[281] = 32'h3ff458cc;
RsqrteLUT[282] = 32'h3ff3e9ca;
RsqrteLUT[283] = 32'h3ff37b5f;
RsqrteLUT[284] = 32'h3ff30d89;
RsqrteLUT[285] = 32'h3ff2a048;
RsqrteLUT[286] = 32'h3ff23399;
RsqrteLUT[287] = 32'h3ff1c77b;
RsqrteLUT[288] = 32'h3ff15bee;
RsqrteLUT[289] = 32'h3ff0f0f0;
RsqrteLUT[290] = 32'h3ff08680;
RsqrteLUT[291] = 32'h3ff01c9d;
RsqrteLUT[292] = 32'h3fefb344;
RsqrteLUT[293] = 32'h3fef4a76;
RsqrteLUT[294] = 32'h3feee231;
RsqrteLUT[295] = 32'h3fee7a74;
RsqrteLUT[296] = 32'h3fee133d;
RsqrteLUT[297] = 32'h3fedac8c;
RsqrteLUT[298] = 32'h3fed4660;
RsqrteLUT[299] = 32'h3fece0b7;
RsqrteLUT[300] = 32'h3fec7b90;
RsqrteLUT[301] = 32'h3fec16ea;
RsqrteLUT[302] = 32'h3febb2c4;
RsqrteLUT[303] = 32'h3feb4f1e;
RsqrteLUT[304] = 32'h3feaebf5;
RsqrteLUT[305] = 32'h3fea8949;
RsqrteLUT[306] = 32'h3fea2719;
RsqrteLUT[307] = 32'h3fe9c564;
RsqrteLUT[308] = 32'h3fe96429;
RsqrteLUT[309] = 32'h3fe90367;
RsqrteLUT[310] = 32'h3fe8a31d;
RsqrteLUT[311] = 32'h3fe8434a;
RsqrteLUT[312] = 32'h3fe7e3ed;
RsqrteLUT[313] = 32'h3fe78505;
RsqrteLUT[314] = 32'h3fe72691;
RsqrteLUT[315] = 32'h3fe6c890;
RsqrteLUT[316] = 32'h3fe66b02;
RsqrteLUT[317] = 32'h3fe60de5;
RsqrteLUT[318] = 32'h3fe5b138;
RsqrteLUT[319] = 32'h3fe554fc;
RsqrteLUT[320] = 32'h3fe4f92e;
RsqrteLUT[321] = 32'h3fe49dce;
RsqrteLUT[322] = 32'h3fe442db;
RsqrteLUT[323] = 32'h3fe3e854;
RsqrteLUT[324] = 32'h3fe38e38;
RsqrteLUT[325] = 32'h3fe33488;
RsqrteLUT[326] = 32'h3fe2db40;
RsqrteLUT[327] = 32'h3fe28262;
RsqrteLUT[328] = 32'h3fe229ec;
RsqrteLUT[329] = 32'h3fe1d1dd;
RsqrteLUT[330] = 32'h3fe17a35;
RsqrteLUT[331] = 32'h3fe122f3;
RsqrteLUT[332] = 32'h3fe0cc15;
RsqrteLUT[333] = 32'h3fe0759c;
RsqrteLUT[334] = 32'h3fe01f86;
RsqrteLUT[335] = 32'h3fdfc9d3;
RsqrteLUT[336] = 32'h3fdf7482;
RsqrteLUT[337] = 32'h3fdf1f93;
RsqrteLUT[338] = 32'h3fdecb03;
RsqrteLUT[339] = 32'h3fde76d4;
RsqrteLUT[340] = 32'h3fde2304;
RsqrteLUT[341] = 32'h3fddcf92;
RsqrteLUT[342] = 32'h3fdd7c7f;
RsqrteLUT[343] = 32'h3fdd29c8;
RsqrteLUT[344] = 32'h3fdcd76d;
RsqrteLUT[345] = 32'h3fdc856f;
RsqrteLUT[346] = 32'h3fdc33cb;
RsqrteLUT[347] = 32'h3fdbe282;
RsqrteLUT[348] = 32'h3fdb9192;
RsqrteLUT[349] = 32'h3fdb40fc;
RsqrteLUT[350] = 32'h3fdaf0be;
RsqrteLUT[351] = 32'h3fdaa0d8;
RsqrteLUT[352] = 32'h3fda5149;
RsqrteLUT[353] = 32'h3fda0211;
RsqrteLUT[354] = 32'h3fd9b32f;
RsqrteLUT[355] = 32'h3fd964a2;
RsqrteLUT[356] = 32'h3fd9166a;
RsqrteLUT[357] = 32'h3fd8c886;
RsqrteLUT[358] = 32'h3fd87af6;
RsqrteLUT[359] = 32'h3fd82db9;
RsqrteLUT[360] = 32'h3fd7e0ce;
RsqrteLUT[361] = 32'h3fd79435;
RsqrteLUT[362] = 32'h3fd747ee;
RsqrteLUT[363] = 32'h3fd6fbf7;
RsqrteLUT[364] = 32'h3fd6b050;
RsqrteLUT[365] = 32'h3fd664f9;
RsqrteLUT[366] = 32'h3fd619f2;
RsqrteLUT[367] = 32'h3fd5cf38;
RsqrteLUT[368] = 32'h3fd584cd;
RsqrteLUT[369] = 32'h3fd53aaf;
RsqrteLUT[370] = 32'h3fd4f0de;
RsqrteLUT[371] = 32'h3fd4a75a;
RsqrteLUT[372] = 32'h3fd45e22;
RsqrteLUT[373] = 32'h3fd41535;
RsqrteLUT[374] = 32'h3fd3cc92;
RsqrteLUT[375] = 32'h3fd3843b;
RsqrteLUT[376] = 32'h3fd33c2d;
RsqrteLUT[377] = 32'h3fd2f469;
RsqrteLUT[378] = 32'h3fd2acee;
RsqrteLUT[379] = 32'h3fd265bb;
RsqrteLUT[380] = 32'h3fd21ed0;
RsqrteLUT[381] = 32'h3fd1d82d;
RsqrteLUT[382] = 32'h3fd191d0;
RsqrteLUT[383] = 32'h3fd14bbb;
RsqrteLUT[384] = 32'h3fd105eb;
RsqrteLUT[385] = 32'h3fd0c061;
RsqrteLUT[386] = 32'h3fd07b1c;
RsqrteLUT[387] = 32'h3fd0361d;
RsqrteLUT[388] = 32'h3fcff161;
RsqrteLUT[389] = 32'h3fcface9;
RsqrteLUT[390] = 32'h3fcf68b5;
RsqrteLUT[391] = 32'h3fcf24c4;
RsqrteLUT[392] = 32'h3fcee115;
RsqrteLUT[393] = 32'h3fce9da9;
RsqrteLUT[394] = 32'h3fce5a7e;
RsqrteLUT[395] = 32'h3fce1795;
RsqrteLUT[396] = 32'h3fcdd4ed;
RsqrteLUT[397] = 32'h3fcd9285;
RsqrteLUT[398] = 32'h3fcd505d;
RsqrteLUT[399] = 32'h3fcd0e75;
RsqrteLUT[400] = 32'h3fcccccc;
RsqrteLUT[401] = 32'h3fcc8b62;
RsqrteLUT[402] = 32'h3fcc4a37;
RsqrteLUT[403] = 32'h3fcc094a;
RsqrteLUT[404] = 32'h3fcbc89b;
RsqrteLUT[405] = 32'h3fcb8829;
RsqrteLUT[406] = 32'h3fcb47f3;
RsqrteLUT[407] = 32'h3fcb07fb;
RsqrteLUT[408] = 32'h3fcac83f;
RsqrteLUT[409] = 32'h3fca88bf;
RsqrteLUT[410] = 32'h3fca497a;
RsqrteLUT[411] = 32'h3fca0a70;
RsqrteLUT[412] = 32'h3fc9cba1;
RsqrteLUT[413] = 32'h3fc98d0d;
RsqrteLUT[414] = 32'h3fc94eb2;
RsqrteLUT[415] = 32'h3fc91092;
RsqrteLUT[416] = 32'h3fc8d2ab;
RsqrteLUT[417] = 32'h3fc894fc;
RsqrteLUT[418] = 32'h3fc85787;
RsqrteLUT[419] = 32'h3fc81a4a;
RsqrteLUT[420] = 32'h3fc7dd45;
RsqrteLUT[421] = 32'h3fc7a077;
RsqrteLUT[422] = 32'h3fc763e1;
RsqrteLUT[423] = 32'h3fc72782;
RsqrteLUT[424] = 32'h3fc6eb5a;
RsqrteLUT[425] = 32'h3fc6af68;
RsqrteLUT[426] = 32'h3fc673ac;
RsqrteLUT[427] = 32'h3fc63826;
RsqrteLUT[428] = 32'h3fc5fcd5;
RsqrteLUT[429] = 32'h3fc5c1b9;
RsqrteLUT[430] = 32'h3fc586d3;
RsqrteLUT[431] = 32'h3fc54c20;
RsqrteLUT[432] = 32'h3fc511a2;
RsqrteLUT[433] = 32'h3fc4d758;
RsqrteLUT[434] = 32'h3fc49d42;
RsqrteLUT[435] = 32'h3fc4635e;
RsqrteLUT[436] = 32'h3fc429ae;
RsqrteLUT[437] = 32'h3fc3f031;
RsqrteLUT[438] = 32'h3fc3b6e6;
RsqrteLUT[439] = 32'h3fc37dcd;
RsqrteLUT[440] = 32'h3fc344e6;
RsqrteLUT[441] = 32'h3fc30c30;
RsqrteLUT[442] = 32'h3fc2d3ac;
RsqrteLUT[443] = 32'h3fc29b59;
RsqrteLUT[444] = 32'h3fc26336;
RsqrteLUT[445] = 32'h3fc22b45;
RsqrteLUT[446] = 32'h3fc1f383;
RsqrteLUT[447] = 32'h3fc1bbf1;
RsqrteLUT[448] = 32'h3fc1848f;
RsqrteLUT[449] = 32'h3fc14d5c;
RsqrteLUT[450] = 32'h3fc11658;
RsqrteLUT[451] = 32'h3fc0df83;
RsqrteLUT[452] = 32'h3fc0a8dd;
RsqrteLUT[453] = 32'h3fc07265;
RsqrteLUT[454] = 32'h3fc03c1c;
RsqrteLUT[455] = 32'h3fc00600;
RsqrteLUT[456] = 32'h3fbfd011;
RsqrteLUT[457] = 32'h3fbf9a51;
RsqrteLUT[458] = 32'h3fbf64bd;
RsqrteLUT[459] = 32'h3fbf2f56;
RsqrteLUT[460] = 32'h3fbefa1b;
RsqrteLUT[461] = 32'h3fbec50d;
RsqrteLUT[462] = 32'h3fbe902b;
RsqrteLUT[463] = 32'h3fbe5b75;
RsqrteLUT[464] = 32'h3fbe26eb;
RsqrteLUT[465] = 32'h3fbdf28c;
RsqrteLUT[466] = 32'h3fbdbe58;
RsqrteLUT[467] = 32'h3fbd8a4f;
RsqrteLUT[468] = 32'h3fbd5671;
RsqrteLUT[469] = 32'h3fbd22bd;
RsqrteLUT[470] = 32'h3fbcef34;
RsqrteLUT[471] = 32'h3fbcbbd4;
RsqrteLUT[472] = 32'h3fbc889f;
RsqrteLUT[473] = 32'h3fbc5593;
RsqrteLUT[474] = 32'h3fbc22b0;
RsqrteLUT[475] = 32'h3fbbeff7;
RsqrteLUT[476] = 32'h3fbbbd66;
RsqrteLUT[477] = 32'h3fbb8aff;
RsqrteLUT[478] = 32'h3fbb58bf;
RsqrteLUT[479] = 32'h3fbb26a9;
RsqrteLUT[480] = 32'h3fbaf4ba;
RsqrteLUT[481] = 32'h3fbac2f3;
RsqrteLUT[482] = 32'h3fba9153;
RsqrteLUT[483] = 32'h3fba5fdc;
RsqrteLUT[484] = 32'h3fba2e8b;
RsqrteLUT[485] = 32'h3fb9fd62;
RsqrteLUT[486] = 32'h3fb9cc5f;
RsqrteLUT[487] = 32'h3fb99b83;
RsqrteLUT[488] = 32'h3fb96ace;
RsqrteLUT[489] = 32'h3fb93a3e;
RsqrteLUT[490] = 32'h3fb909d5;
RsqrteLUT[491] = 32'h3fb8d992;
RsqrteLUT[492] = 32'h3fb8a974;
RsqrteLUT[493] = 32'h3fb8797c;
RsqrteLUT[494] = 32'h3fb849aa;
RsqrteLUT[495] = 32'h3fb819fc;
RsqrteLUT[496] = 32'h3fb7ea73;
RsqrteLUT[497] = 32'h3fb7bb0f;
RsqrteLUT[498] = 32'h3fb78bd0;
RsqrteLUT[499] = 32'h3fb75cb5;
RsqrteLUT[500] = 32'h3fb72dbe;
RsqrteLUT[501] = 32'h3fb6feeb;
RsqrteLUT[502] = 32'h3fb6d03c;
RsqrteLUT[503] = 32'h3fb6a1b1;
RsqrteLUT[504] = 32'h3fb67349;
RsqrteLUT[505] = 32'h3fb64505;
RsqrteLUT[506] = 32'h3fb616e3;
RsqrteLUT[507] = 32'h3fb5e8e5;
RsqrteLUT[508] = 32'h3fb5bb09;
RsqrteLUT[509] = 32'h3fb58d50;
RsqrteLUT[510] = 32'h3fb55fb9;
RsqrteLUT[511] = 32'h3fb53245;
RsqrteLUT[512] = 32'h3fb504f3;
RsqrteLUT[513] = 32'h3fb4d7c2;
RsqrteLUT[514] = 32'h3fb4aab4;
RsqrteLUT[515] = 32'h3fb47dc7;
RsqrteLUT[516] = 32'h3fb450fc;
RsqrteLUT[517] = 32'h3fb42451;
RsqrteLUT[518] = 32'h3fb3f7c8;
RsqrteLUT[519] = 32'h3fb3cb60;
RsqrteLUT[520] = 32'h3fb39f19;
RsqrteLUT[521] = 32'h3fb372f2;
RsqrteLUT[522] = 32'h3fb346ec;
RsqrteLUT[523] = 32'h3fb31b06;
RsqrteLUT[524] = 32'h3fb2ef41;
RsqrteLUT[525] = 32'h3fb2c39b;
RsqrteLUT[526] = 32'h3fb29816;
RsqrteLUT[527] = 32'h3fb26cb0;
RsqrteLUT[528] = 32'h3fb24169;
RsqrteLUT[529] = 32'h3fb21642;
RsqrteLUT[530] = 32'h3fb1eb3b;
RsqrteLUT[531] = 32'h3fb1c052;
RsqrteLUT[532] = 32'h3fb19589;
RsqrteLUT[533] = 32'h3fb16ade;
RsqrteLUT[534] = 32'h3fb14052;
RsqrteLUT[535] = 32'h3fb115e4;
RsqrteLUT[536] = 32'h3fb0eb95;
RsqrteLUT[537] = 32'h3fb0c164;
RsqrteLUT[538] = 32'h3fb09752;
RsqrteLUT[539] = 32'h3fb06d5d;
RsqrteLUT[540] = 32'h3fb04386;
RsqrteLUT[541] = 32'h3fb019cd;
RsqrteLUT[542] = 32'h3faff032;
RsqrteLUT[543] = 32'h3fafc6b4;
RsqrteLUT[544] = 32'h3faf9d53;
RsqrteLUT[545] = 32'h3faf740f;
RsqrteLUT[546] = 32'h3faf4ae8;
RsqrteLUT[547] = 32'h3faf21df;
RsqrteLUT[548] = 32'h3faef8f2;
RsqrteLUT[549] = 32'h3faed022;
RsqrteLUT[550] = 32'h3faea76e;
RsqrteLUT[551] = 32'h3fae7ed6;
RsqrteLUT[552] = 32'h3fae565b;
RsqrteLUT[553] = 32'h3fae2dfc;
RsqrteLUT[554] = 32'h3fae05b9;
RsqrteLUT[555] = 32'h3faddd92;
RsqrteLUT[556] = 32'h3fadb587;
RsqrteLUT[557] = 32'h3fad8d97;
RsqrteLUT[558] = 32'h3fad65c3;
RsqrteLUT[559] = 32'h3fad3e0a;
RsqrteLUT[560] = 32'h3fad166c;
RsqrteLUT[561] = 32'h3faceee9;
RsqrteLUT[562] = 32'h3facc782;
RsqrteLUT[563] = 32'h3faca035;
RsqrteLUT[564] = 32'h3fac7903;
RsqrteLUT[565] = 32'h3fac51ec;
RsqrteLUT[566] = 32'h3fac2aef;
RsqrteLUT[567] = 32'h3fac040d;
RsqrteLUT[568] = 32'h3fabdd45;
RsqrteLUT[569] = 32'h3fabb697;
RsqrteLUT[570] = 32'h3fab9003;
RsqrteLUT[571] = 32'h3fab698a;
RsqrteLUT[572] = 32'h3fab432a;
RsqrteLUT[573] = 32'h3fab1ce4;
RsqrteLUT[574] = 32'h3faaf6b7;
RsqrteLUT[575] = 32'h3faad0a4;
RsqrteLUT[576] = 32'h3faaaaaa;
RsqrteLUT[577] = 32'h3faa84ca;
RsqrteLUT[578] = 32'h3faa5f03;
RsqrteLUT[579] = 32'h3faa3954;
RsqrteLUT[580] = 32'h3faa13bf;
RsqrteLUT[581] = 32'h3fa9ee43;
RsqrteLUT[582] = 32'h3fa9c8df;
RsqrteLUT[583] = 32'h3fa9a394;
RsqrteLUT[584] = 32'h3fa97e62;
RsqrteLUT[585] = 32'h3fa95948;
RsqrteLUT[586] = 32'h3fa93446;
RsqrteLUT[587] = 32'h3fa90f5c;
RsqrteLUT[588] = 32'h3fa8ea8b;
RsqrteLUT[589] = 32'h3fa8c5d2;
RsqrteLUT[590] = 32'h3fa8a130;
RsqrteLUT[591] = 32'h3fa87ca7;
RsqrteLUT[592] = 32'h3fa85835;
RsqrteLUT[593] = 32'h3fa833da;
RsqrteLUT[594] = 32'h3fa80f98;
RsqrteLUT[595] = 32'h3fa7eb6c;
RsqrteLUT[596] = 32'h3fa7c758;
RsqrteLUT[597] = 32'h3fa7a35b;
RsqrteLUT[598] = 32'h3fa77f76;
RsqrteLUT[599] = 32'h3fa75ba7;
RsqrteLUT[600] = 32'h3fa737ef;
RsqrteLUT[601] = 32'h3fa7144e;
RsqrteLUT[602] = 32'h3fa6f0c4;
RsqrteLUT[603] = 32'h3fa6cd50;
RsqrteLUT[604] = 32'h3fa6a9f3;
RsqrteLUT[605] = 32'h3fa686ad;
RsqrteLUT[606] = 32'h3fa6637d;
RsqrteLUT[607] = 32'h3fa64063;
RsqrteLUT[608] = 32'h3fa61d5f;
RsqrteLUT[609] = 32'h3fa5fa71;
RsqrteLUT[610] = 32'h3fa5d799;
RsqrteLUT[611] = 32'h3fa5b4d8;
RsqrteLUT[612] = 32'h3fa5922c;
RsqrteLUT[613] = 32'h3fa56f95;
RsqrteLUT[614] = 32'h3fa54d15;
RsqrteLUT[615] = 32'h3fa52aaa;
RsqrteLUT[616] = 32'h3fa50854;
RsqrteLUT[617] = 32'h3fa4e614;
RsqrteLUT[618] = 32'h3fa4c3e9;
RsqrteLUT[619] = 32'h3fa4a1d3;
RsqrteLUT[620] = 32'h3fa47fd3;
RsqrteLUT[621] = 32'h3fa45de7;
RsqrteLUT[622] = 32'h3fa43c11;
RsqrteLUT[623] = 32'h3fa41a4f;
RsqrteLUT[624] = 32'h3fa3f8a2;
RsqrteLUT[625] = 32'h3fa3d70a;
RsqrteLUT[626] = 32'h3fa3b586;
RsqrteLUT[627] = 32'h3fa39417;
RsqrteLUT[628] = 32'h3fa372bc;
RsqrteLUT[629] = 32'h3fa35176;
RsqrteLUT[630] = 32'h3fa33044;
RsqrteLUT[631] = 32'h3fa30f26;
RsqrteLUT[632] = 32'h3fa2ee1d;
RsqrteLUT[633] = 32'h3fa2cd27;
RsqrteLUT[634] = 32'h3fa2ac45;
RsqrteLUT[635] = 32'h3fa28b78;
RsqrteLUT[636] = 32'h3fa26abe;
RsqrteLUT[637] = 32'h3fa24a18;
RsqrteLUT[638] = 32'h3fa22985;
RsqrteLUT[639] = 32'h3fa20906;
RsqrteLUT[640] = 32'h3fa1e89b;
RsqrteLUT[641] = 32'h3fa1c843;
RsqrteLUT[642] = 32'h3fa1a7fe;
RsqrteLUT[643] = 32'h3fa187cc;
RsqrteLUT[644] = 32'h3fa167ae;
RsqrteLUT[645] = 32'h3fa147a3;
RsqrteLUT[646] = 32'h3fa127ab;
RsqrteLUT[647] = 32'h3fa107c6;
RsqrteLUT[648] = 32'h3fa0e7f4;
RsqrteLUT[649] = 32'h3fa0c835;
RsqrteLUT[650] = 32'h3fa0a888;
RsqrteLUT[651] = 32'h3fa088ef;
RsqrteLUT[652] = 32'h3fa06967;
RsqrteLUT[653] = 32'h3fa049f3;
RsqrteLUT[654] = 32'h3fa02a90;
RsqrteLUT[655] = 32'h3fa00b41;
RsqrteLUT[656] = 32'h3f9fec03;
RsqrteLUT[657] = 32'h3f9fccd8;
RsqrteLUT[658] = 32'h3f9fadbf;
RsqrteLUT[659] = 32'h3f9f8eb8;
RsqrteLUT[660] = 32'h3f9f6fc3;
RsqrteLUT[661] = 32'h3f9f50e1;
RsqrteLUT[662] = 32'h3f9f3210;
RsqrteLUT[663] = 32'h3f9f1351;
RsqrteLUT[664] = 32'h3f9ef4a4;
RsqrteLUT[665] = 32'h3f9ed608;
RsqrteLUT[666] = 32'h3f9eb77e;
RsqrteLUT[667] = 32'h3f9e9906;
RsqrteLUT[668] = 32'h3f9e7a9f;
RsqrteLUT[669] = 32'h3f9e5c4a;
RsqrteLUT[670] = 32'h3f9e3e06;
RsqrteLUT[671] = 32'h3f9e1fd3;
RsqrteLUT[672] = 32'h3f9e01b2;
RsqrteLUT[673] = 32'h3f9de3a2;
RsqrteLUT[674] = 32'h3f9dc5a3;
RsqrteLUT[675] = 32'h3f9da7b5;
RsqrteLUT[676] = 32'h3f9d89d8;
RsqrteLUT[677] = 32'h3f9d6c0c;
RsqrteLUT[678] = 32'h3f9d4e51;
RsqrteLUT[679] = 32'h3f9d30a7;
RsqrteLUT[680] = 32'h3f9d130d;
RsqrteLUT[681] = 32'h3f9cf585;
RsqrteLUT[682] = 32'h3f9cd80c;
RsqrteLUT[683] = 32'h3f9cbaa5;
RsqrteLUT[684] = 32'h3f9c9d4e;
RsqrteLUT[685] = 32'h3f9c8007;
RsqrteLUT[686] = 32'h3f9c62d1;
RsqrteLUT[687] = 32'h3f9c45ab;
RsqrteLUT[688] = 32'h3f9c2895;
RsqrteLUT[689] = 32'h3f9c0b90;
RsqrteLUT[690] = 32'h3f9bee9b;
RsqrteLUT[691] = 32'h3f9bd1b6;
RsqrteLUT[692] = 32'h3f9bb4e0;
RsqrteLUT[693] = 32'h3f9b981b;
RsqrteLUT[694] = 32'h3f9b7b66;
RsqrteLUT[695] = 32'h3f9b5ec1;
RsqrteLUT[696] = 32'h3f9b422b;
RsqrteLUT[697] = 32'h3f9b25a5;
RsqrteLUT[698] = 32'h3f9b092f;
RsqrteLUT[699] = 32'h3f9aecc9;
RsqrteLUT[700] = 32'h3f9ad072;
RsqrteLUT[701] = 32'h3f9ab42b;
RsqrteLUT[702] = 32'h3f9a97f3;
RsqrteLUT[703] = 32'h3f9a7bca;
RsqrteLUT[704] = 32'h3f9a5fb1;
RsqrteLUT[705] = 32'h3f9a43a8;
RsqrteLUT[706] = 32'h3f9a27ad;
RsqrteLUT[707] = 32'h3f9a0bc2;
RsqrteLUT[708] = 32'h3f99efe6;
RsqrteLUT[709] = 32'h3f99d419;
RsqrteLUT[710] = 32'h3f99b85b;
RsqrteLUT[711] = 32'h3f999cac;
RsqrteLUT[712] = 32'h3f99810c;
RsqrteLUT[713] = 32'h3f99657a;
RsqrteLUT[714] = 32'h3f9949f8;
RsqrteLUT[715] = 32'h3f992e84;
RsqrteLUT[716] = 32'h3f99131f;
RsqrteLUT[717] = 32'h3f98f7c9;
RsqrteLUT[718] = 32'h3f98dc82;
RsqrteLUT[719] = 32'h3f98c149;
RsqrteLUT[720] = 32'h3f98a61e;
RsqrteLUT[721] = 32'h3f988b02;
RsqrteLUT[722] = 32'h3f986ff5;
RsqrteLUT[723] = 32'h3f9854f6;
RsqrteLUT[724] = 32'h3f983a05;
RsqrteLUT[725] = 32'h3f981f22;
RsqrteLUT[726] = 32'h3f98044e;
RsqrteLUT[727] = 32'h3f97e987;
RsqrteLUT[728] = 32'h3f97cecf;
RsqrteLUT[729] = 32'h3f97b425;
RsqrteLUT[730] = 32'h3f979989;
RsqrteLUT[731] = 32'h3f977efb;
RsqrteLUT[732] = 32'h3f97647b;
RsqrteLUT[733] = 32'h3f974a09;
RsqrteLUT[734] = 32'h3f972fa5;
RsqrteLUT[735] = 32'h3f97154e;
RsqrteLUT[736] = 32'h3f96fb06;
RsqrteLUT[737] = 32'h3f96e0cb;
RsqrteLUT[738] = 32'h3f96c69d;
RsqrteLUT[739] = 32'h3f96ac7d;
RsqrteLUT[740] = 32'h3f96926b;
RsqrteLUT[741] = 32'h3f967866;
RsqrteLUT[742] = 32'h3f965e6f;
RsqrteLUT[743] = 32'h3f964485;
RsqrteLUT[744] = 32'h3f962aa9;
RsqrteLUT[745] = 32'h3f9610da;
RsqrteLUT[746] = 32'h3f95f718;
RsqrteLUT[747] = 32'h3f95dd63;
RsqrteLUT[748] = 32'h3f95c3bc;
RsqrteLUT[749] = 32'h3f95aa22;
RsqrteLUT[750] = 32'h3f959094;
RsqrteLUT[751] = 32'h3f957714;
RsqrteLUT[752] = 32'h3f955da1;
RsqrteLUT[753] = 32'h3f95443b;
RsqrteLUT[754] = 32'h3f952ae2;
RsqrteLUT[755] = 32'h3f951196;
RsqrteLUT[756] = 32'h3f94f857;
RsqrteLUT[757] = 32'h3f94df24;
RsqrteLUT[758] = 32'h3f94c5fe;
RsqrteLUT[759] = 32'h3f94ace5;
RsqrteLUT[760] = 32'h3f9493d9;
RsqrteLUT[761] = 32'h3f947ad9;
RsqrteLUT[762] = 32'h3f9461e6;
RsqrteLUT[763] = 32'h3f9448ff;
RsqrteLUT[764] = 32'h3f943025;
RsqrteLUT[765] = 32'h3f941758;
RsqrteLUT[766] = 32'h3f93fe97;
RsqrteLUT[767] = 32'h3f93e5e2;
RsqrteLUT[768] = 32'h3f93cd3a;
RsqrteLUT[769] = 32'h3f93b49e;
RsqrteLUT[770] = 32'h3f939c0e;
RsqrteLUT[771] = 32'h3f93838a;
RsqrteLUT[772] = 32'h3f936b13;
RsqrteLUT[773] = 32'h3f9352a8;
RsqrteLUT[774] = 32'h3f933a49;
RsqrteLUT[775] = 32'h3f9321f6;
RsqrteLUT[776] = 32'h3f9309af;
RsqrteLUT[777] = 32'h3f92f174;
RsqrteLUT[778] = 32'h3f92d945;
RsqrteLUT[779] = 32'h3f92c122;
RsqrteLUT[780] = 32'h3f92a90b;
RsqrteLUT[781] = 32'h3f9290ff;
RsqrteLUT[782] = 32'h3f927900;
RsqrteLUT[783] = 32'h3f92610c;
RsqrteLUT[784] = 32'h3f924924;
RsqrteLUT[785] = 32'h3f923148;
RsqrteLUT[786] = 32'h3f921977;
RsqrteLUT[787] = 32'h3f9201b2;
RsqrteLUT[788] = 32'h3f91e9f9;
RsqrteLUT[789] = 32'h3f91d24b;
RsqrteLUT[790] = 32'h3f91baa8;
RsqrteLUT[791] = 32'h3f91a312;
RsqrteLUT[792] = 32'h3f918b86;
RsqrteLUT[793] = 32'h3f917406;
RsqrteLUT[794] = 32'h3f915c91;
RsqrteLUT[795] = 32'h3f914528;
RsqrteLUT[796] = 32'h3f912dca;
RsqrteLUT[797] = 32'h3f911677;
RsqrteLUT[798] = 32'h3f90ff30;
RsqrteLUT[799] = 32'h3f90e7f3;
RsqrteLUT[800] = 32'h3f90d0c2;
RsqrteLUT[801] = 32'h3f90b99c;
RsqrteLUT[802] = 32'h3f90a281;
RsqrteLUT[803] = 32'h3f908b71;
RsqrteLUT[804] = 32'h3f90746c;
RsqrteLUT[805] = 32'h3f905d72;
RsqrteLUT[806] = 32'h3f904683;
RsqrteLUT[807] = 32'h3f902f9f;
RsqrteLUT[808] = 32'h3f9018c6;
RsqrteLUT[809] = 32'h3f9001f8;
RsqrteLUT[810] = 32'h3f8feb34;
RsqrteLUT[811] = 32'h3f8fd47b;
RsqrteLUT[812] = 32'h3f8fbdcd;
RsqrteLUT[813] = 32'h3f8fa72a;
RsqrteLUT[814] = 32'h3f8f9091;
RsqrteLUT[815] = 32'h3f8f7a03;
RsqrteLUT[816] = 32'h3f8f6380;
RsqrteLUT[817] = 32'h3f8f4d07;
RsqrteLUT[818] = 32'h3f8f3699;
RsqrteLUT[819] = 32'h3f8f2035;
RsqrteLUT[820] = 32'h3f8f09dc;
RsqrteLUT[821] = 32'h3f8ef38e;
RsqrteLUT[822] = 32'h3f8edd49;
RsqrteLUT[823] = 32'h3f8ec70f;
RsqrteLUT[824] = 32'h3f8eb0e0;
RsqrteLUT[825] = 32'h3f8e9aba;
RsqrteLUT[826] = 32'h3f8e84a0;
RsqrteLUT[827] = 32'h3f8e6e8f;
RsqrteLUT[828] = 32'h3f8e5888;
RsqrteLUT[829] = 32'h3f8e428c;
RsqrteLUT[830] = 32'h3f8e2c9a;
RsqrteLUT[831] = 32'h3f8e16b2;
RsqrteLUT[832] = 32'h3f8e00d5;
RsqrteLUT[833] = 32'h3f8deb01;
RsqrteLUT[834] = 32'h3f8dd537;
RsqrteLUT[835] = 32'h3f8dbf78;
RsqrteLUT[836] = 32'h3f8da9c2;
RsqrteLUT[837] = 32'h3f8d9416;
RsqrteLUT[838] = 32'h3f8d7e74;
RsqrteLUT[839] = 32'h3f8d68dd;
RsqrteLUT[840] = 32'h3f8d534f;
RsqrteLUT[841] = 32'h3f8d3dcb;
RsqrteLUT[842] = 32'h3f8d2850;
RsqrteLUT[843] = 32'h3f8d12e0;
RsqrteLUT[844] = 32'h3f8cfd79;
RsqrteLUT[845] = 32'h3f8ce81c;
RsqrteLUT[846] = 32'h3f8cd2c9;
RsqrteLUT[847] = 32'h3f8cbd7f;
RsqrteLUT[848] = 32'h3f8ca83f;
RsqrteLUT[849] = 32'h3f8c9309;
RsqrteLUT[850] = 32'h3f8c7ddc;
RsqrteLUT[851] = 32'h3f8c68b8;
RsqrteLUT[852] = 32'h3f8c539f;
RsqrteLUT[853] = 32'h3f8c3e8e;
RsqrteLUT[854] = 32'h3f8c2988;
RsqrteLUT[855] = 32'h3f8c148a;
RsqrteLUT[856] = 32'h3f8bff97;
RsqrteLUT[857] = 32'h3f8beaac;
RsqrteLUT[858] = 32'h3f8bd5cb;
RsqrteLUT[859] = 32'h3f8bc0f3;
RsqrteLUT[860] = 32'h3f8bac25;
RsqrteLUT[861] = 32'h3f8b975f;
RsqrteLUT[862] = 32'h3f8b82a3;
RsqrteLUT[863] = 32'h3f8b6df1;
RsqrteLUT[864] = 32'h3f8b5947;
RsqrteLUT[865] = 32'h3f8b44a7;
RsqrteLUT[866] = 32'h3f8b3010;
RsqrteLUT[867] = 32'h3f8b1b82;
RsqrteLUT[868] = 32'h3f8b06fd;
RsqrteLUT[869] = 32'h3f8af281;
RsqrteLUT[870] = 32'h3f8ade0e;
RsqrteLUT[871] = 32'h3f8ac9a4;
RsqrteLUT[872] = 32'h3f8ab543;
RsqrteLUT[873] = 32'h3f8aa0eb;
RsqrteLUT[874] = 32'h3f8a8c9c;
RsqrteLUT[875] = 32'h3f8a7856;
RsqrteLUT[876] = 32'h3f8a6419;
RsqrteLUT[877] = 32'h3f8a4fe5;
RsqrteLUT[878] = 32'h3f8a3bb9;
RsqrteLUT[879] = 32'h3f8a2797;
RsqrteLUT[880] = 32'h3f8a137d;
RsqrteLUT[881] = 32'h3f89ff6c;
RsqrteLUT[882] = 32'h3f89eb63;
RsqrteLUT[883] = 32'h3f89d764;
RsqrteLUT[884] = 32'h3f89c36d;
RsqrteLUT[885] = 32'h3f89af7f;
RsqrteLUT[886] = 32'h3f899b99;
RsqrteLUT[887] = 32'h3f8987bc;
RsqrteLUT[888] = 32'h3f8973e8;
RsqrteLUT[889] = 32'h3f89601c;
RsqrteLUT[890] = 32'h3f894c58;
RsqrteLUT[891] = 32'h3f89389e;
RsqrteLUT[892] = 32'h3f8924eb;
RsqrteLUT[893] = 32'h3f891142;
RsqrteLUT[894] = 32'h3f88fda0;
RsqrteLUT[895] = 32'h3f88ea07;
RsqrteLUT[896] = 32'h3f88d677;
RsqrteLUT[897] = 32'h3f88c2ef;
RsqrteLUT[898] = 32'h3f88af6f;
RsqrteLUT[899] = 32'h3f889bf7;
RsqrteLUT[900] = 32'h3f888888;
RsqrteLUT[901] = 32'h3f887521;
RsqrteLUT[902] = 32'h3f8861c3;
RsqrteLUT[903] = 32'h3f884e6c;
RsqrteLUT[904] = 32'h3f883b1e;
RsqrteLUT[905] = 32'h3f8827d8;
RsqrteLUT[906] = 32'h3f88149a;
RsqrteLUT[907] = 32'h3f880165;
RsqrteLUT[908] = 32'h3f87ee37;
RsqrteLUT[909] = 32'h3f87db12;
RsqrteLUT[910] = 32'h3f87c7f4;
RsqrteLUT[911] = 32'h3f87b4df;
RsqrteLUT[912] = 32'h3f87a1d2;
RsqrteLUT[913] = 32'h3f878ecc;
RsqrteLUT[914] = 32'h3f877bcf;
RsqrteLUT[915] = 32'h3f8768da;
RsqrteLUT[916] = 32'h3f8755ed;
RsqrteLUT[917] = 32'h3f874307;
RsqrteLUT[918] = 32'h3f87302a;
RsqrteLUT[919] = 32'h3f871d54;
RsqrteLUT[920] = 32'h3f870a86;
RsqrteLUT[921] = 32'h3f86f7c1;
RsqrteLUT[922] = 32'h3f86e502;
RsqrteLUT[923] = 32'h3f86d24c;
RsqrteLUT[924] = 32'h3f86bf9e;
RsqrteLUT[925] = 32'h3f86acf7;
RsqrteLUT[926] = 32'h3f869a58;
RsqrteLUT[927] = 32'h3f8687c1;
RsqrteLUT[928] = 32'h3f867531;
RsqrteLUT[929] = 32'h3f8662a9;
RsqrteLUT[930] = 32'h3f865029;
RsqrteLUT[931] = 32'h3f863db0;
RsqrteLUT[932] = 32'h3f862b3f;
RsqrteLUT[933] = 32'h3f8618d6;
RsqrteLUT[934] = 32'h3f860674;
RsqrteLUT[935] = 32'h3f85f41a;
RsqrteLUT[936] = 32'h3f85e1c7;
RsqrteLUT[937] = 32'h3f85cf7c;
RsqrteLUT[938] = 32'h3f85bd38;
RsqrteLUT[939] = 32'h3f85aafc;
RsqrteLUT[940] = 32'h3f8598c7;
RsqrteLUT[941] = 32'h3f858699;
RsqrteLUT[942] = 32'h3f857473;
RsqrteLUT[943] = 32'h3f856255;
RsqrteLUT[944] = 32'h3f85503d;
RsqrteLUT[945] = 32'h3f853e2e;
RsqrteLUT[946] = 32'h3f852c25;
RsqrteLUT[947] = 32'h3f851a24;
RsqrteLUT[948] = 32'h3f85082a;
RsqrteLUT[949] = 32'h3f84f637;
RsqrteLUT[950] = 32'h3f84e44c;
RsqrteLUT[951] = 32'h3f84d268;
RsqrteLUT[952] = 32'h3f84c08b;
RsqrteLUT[953] = 32'h3f84aeb5;
RsqrteLUT[954] = 32'h3f849ce6;
RsqrteLUT[955] = 32'h3f848b1f;
RsqrteLUT[956] = 32'h3f84795f;
RsqrteLUT[957] = 32'h3f8467a5;
RsqrteLUT[958] = 32'h3f8455f3;
RsqrteLUT[959] = 32'h3f844448;
RsqrteLUT[960] = 32'h3f8432a5;
RsqrteLUT[961] = 32'h3f842108;
RsqrteLUT[962] = 32'h3f840f72;
RsqrteLUT[963] = 32'h3f83fde3;
RsqrteLUT[964] = 32'h3f83ec5b;
RsqrteLUT[965] = 32'h3f83dadb;
RsqrteLUT[966] = 32'h3f83c961;
RsqrteLUT[967] = 32'h3f83b7ee;
RsqrteLUT[968] = 32'h3f83a682;
RsqrteLUT[969] = 32'h3f83951d;
RsqrteLUT[970] = 32'h3f8383bf;
RsqrteLUT[971] = 32'h3f837267;
RsqrteLUT[972] = 32'h3f836117;
RsqrteLUT[973] = 32'h3f834fcd;
RsqrteLUT[974] = 32'h3f833e8a;
RsqrteLUT[975] = 32'h3f832d4e;
RsqrteLUT[976] = 32'h3f831c19;
RsqrteLUT[977] = 32'h3f830aeb;
RsqrteLUT[978] = 32'h3f82f9c3;
RsqrteLUT[979] = 32'h3f82e8a2;
RsqrteLUT[980] = 32'h3f82d788;
RsqrteLUT[981] = 32'h3f82c674;
RsqrteLUT[982] = 32'h3f82b567;
RsqrteLUT[983] = 32'h3f82a461;
RsqrteLUT[984] = 32'h3f829361;
RsqrteLUT[985] = 32'h3f828268;
RsqrteLUT[986] = 32'h3f827176;
RsqrteLUT[987] = 32'h3f82608a;
RsqrteLUT[988] = 32'h3f824fa5;
RsqrteLUT[989] = 32'h3f823ec6;
RsqrteLUT[990] = 32'h3f822dee;
RsqrteLUT[991] = 32'h3f821d1d;
RsqrteLUT[992] = 32'h3f820c52;
RsqrteLUT[993] = 32'h3f81fb8d;
RsqrteLUT[994] = 32'h3f81eacf;
RsqrteLUT[995] = 32'h3f81da18;
RsqrteLUT[996] = 32'h3f81c966;
RsqrteLUT[997] = 32'h3f81b8bc;
RsqrteLUT[998] = 32'h3f81a817;
RsqrteLUT[999] = 32'h3f819779;
RsqrteLUT[1000] = 32'h3f8186e2;
RsqrteLUT[1001] = 32'h3f817651;
RsqrteLUT[1002] = 32'h3f8165c6;
RsqrteLUT[1003] = 32'h3f815542;
RsqrteLUT[1004] = 32'h3f8144c3;
RsqrteLUT[1005] = 32'h3f81344c;
RsqrteLUT[1006] = 32'h3f8123da;
RsqrteLUT[1007] = 32'h3f81136f;
RsqrteLUT[1008] = 32'h3f81030a;
RsqrteLUT[1009] = 32'h3f80f2ab;
RsqrteLUT[1010] = 32'h3f80e252;
RsqrteLUT[1011] = 32'h3f80d200;
RsqrteLUT[1012] = 32'h3f80c1b4;
RsqrteLUT[1013] = 32'h3f80b16e;
RsqrteLUT[1014] = 32'h3f80a12e;
RsqrteLUT[1015] = 32'h3f8090f4;
RsqrteLUT[1016] = 32'h3f8080c1;
RsqrteLUT[1017] = 32'h3f807093;
RsqrteLUT[1018] = 32'h3f80606c;
RsqrteLUT[1019] = 32'h3f80504b;
RsqrteLUT[1020] = 32'h3f804030;
RsqrteLUT[1021] = 32'h3f80301b;
RsqrteLUT[1022] = 32'h3f80200c;
RsqrteLUT[1023] = 32'h3f801003;