
package rf6809_pkg;

typedef logic [23:0] Address;
typedef logic [11:0] Data;

parameter bitsPerByte =	$bits(Data);
parameter BPB = bitsPerByte;
parameter BPBM1 =	BPB-1;
parameter BPBX2M1 =	BPB*2-1;

// The following allows asynchronous reads for icache updating.
// It increases the size of the core.
//`define SUPPORT_AREAD	1

// The following includes an instruction buffer when icache is
// not used.
//`define SUPPORT_IBUF	1

// The following enables support for the checkpoint interrupt.
//`define SUPPORT_CHECKPOINT

//`define EIGHTBIT	1
`define TWELVEBIT	2

`ifdef EIGHTBIT
`define LOBYTE	7:0
`define HIBYTE	15:8
`define DBLBYTE	15:0
`define TRPBYTE		23:0
`define BYTE1		7:0
`define BYTE2		15:8
`define BYTE3		23:16
`define BYTE4		31:24
`define BYTE5		39:32
`define QUINBYTE	47:0
`define HEXBYTE		55:0
`define DBLBYTEP1	16:0
`define LOBYTEP1	8:0
`define HCBIT		3
`endif

`ifdef TWELVEBIT
`define LOBYTE	11:0
`define HIBYTE	23:12
`define DBLBYTE	23:0
`define TRPBYTE		35:0
`define BYTE1		11:0
`define BYTE2		23:12
`define BYTE3		35:24
`define BYTE4		47:36
`define BYTE5		59:48
`define QUINBYTE	59:0
`define HEXBYTE		71:0
`define DBLBYTEP1	24:0
`define LOBYTEP1	12:0
`define HCBIT		3
`endif

`define TRUE		1'b1
`define FALSE		1'b0

`define RST_VECT	24'hFFFFFE
`define NMI_VECT	24'hFFFFFC
`define SWI_VECT	24'hFFFFFA
`define IRQ_VECT	24'hFFFFF8
`define FIRQ_VECT	24'hFFFFF6
`define SWI2_VECT	24'hFFFFF4
`define SWI3_VECT	24'hFFFFF2
`define RESV_VECT	24'hFFFFF0

`define NEG_DP		12'h000
`define OIM_DP		12'h001
`define AIM_DP		12'h002
`define COM_DP		12'h003
`define LSR_DP		12'h004
`define EIM_DP		12'h005
`define ROR_DP		12'h006
`define ASR_DP		12'h007
`define ASL_DP		12'h008
`define ROL_DP		12'h009
`define DEC_DP		12'h00A
`define TIM_DP		12'h00B
`define INC_DP		12'h00C
`define TST_DP		12'h00D
`define JMP_DP		12'h00E
`define CLR_DP		12'h00F

`define PG2			12'h010
`define PG3			12'h011
`define NOP			12'h012
`define SYNC		12'h013
`define SEXW		12'h014
`define FAR			12'h015
`define LBRA		12'h016
`define LBSR		12'h017
`define DAA			12'h019
`define ORCC		12'h01A
`define OUTER		12'h01B
`define ANDCC		12'h01C
`define SEX			12'h01D
`define EXG			12'h01E
`define TFR			12'h01F

`define BRA			12'h020
`define BRN			12'h021
`define BHI			12'h022
`define BLS			12'h023
`define BHS			12'h024
`define BLO			12'h025
`define BNE			12'h026
`define BEQ			12'h027
`define BVC			12'h028
`define BVS			12'h029
`define BPL			12'h02A
`define BMI			12'h02B
`define BGE			12'h02C
`define BLT			12'h02D
`define BGT			12'h02E
`define BLE			12'h02F

`define LEAX_NDX	12'h030
`define LEAY_NDX	12'h031
`define LEAS_NDX	12'h032
`define LEAU_NDX	12'h033
`define PSHS		12'h034
`define PULS		12'h035
`define PSHU		12'h036
`define PULU		12'h037
`define RTF			12'h038
`define RTS			12'h039
`define ABX			12'h03A
`define RTI			12'h03B
`define CWAI		12'h03C
`define MUL			12'h03D
`define SWI			12'h03F

`define NEGA		12'h040
`define COMA		12'h043
`define LSRA		12'h044
`define RORA		12'h046
`define ASRA		12'h047
`define ASLA		12'h048
`define ROLA		12'h049
`define DECA		12'h04A
`define INCA		12'h04C
`define TSTA		12'h04D
`define CLRA		12'h04F

`define NEGB		12'h050
`define COMB		12'h053
`define LSRB		12'h054
`define RORB		12'h056
`define ASRB		12'h057
`define ASLB		12'h058
`define ROLB		12'h059
`define DECB		12'h05A
`define INCB		12'h05C
`define TSTB		12'h05D
`define CLRB		12'h05F

`define NEG_NDX		12'h060
`define OIM_NDX		12'h061
`define AIM_NDX		12'h062
`define COM_NDX		12'h063
`define LSR_NDX		12'h064
`define EIM_NDX		12'h065
`define ROR_NDX		12'h066
`define ASR_NDX		12'h067
`define ASL_NDX		12'h068
`define ROL_NDX		12'h069
`define DEC_NDX		12'h06A
`define TIM_NDX		12'h06B
`define INC_NDX		12'h06C
`define TST_NDX		12'h06D
`define JMP_NDX		12'h06E
`define CLR_NDX		12'h06F

`define NEG_EXT		12'h070
`define OIM_EXT		12'h071
`define AIM_EXT		12'h072
`define COM_EXT		12'h073
`define LSR_EXT		12'h074
`define EIM_EXT		12'h075
`define ROR_EXT		12'h076
`define ASR_EXT		12'h077
`define ASL_EXT		12'h078
`define ROL_EXT		12'h079
`define DEC_EXT		12'h07A
`define TIM_EXT		12'h07B
`define INC_EXT		12'h07C
`define TST_EXT		12'h07D
`define JMP_EXT		12'h07E
`define CLR_EXT		12'h07F

`define SUBA_IMM	12'h080
`define CMPA_IMM	12'h081
`define SBCA_IMM	12'h082
`define SUBD_IMM	12'h083
`define ANDA_IMM	12'h084
`define BITA_IMM	12'h085
`define LDA_IMM		12'h086
`define EORA_IMM	12'h088
`define ADCA_IMM	12'h089
`define ORA_IMM		12'h08A
`define ADDA_IMM	12'h08B
`define CMPX_IMM	12'h08C
`define BSR			12'h08D
`define LDX_IMM		12'h08E
`define JMP_FAR		12'h08F

`define SUBA_DP		12'h090
`define CMPA_DP		12'h091
`define SBCA_DP		12'h092
`define SUBD_DP		12'h093
`define ANDA_DP		12'h094
`define BITA_DP		12'h095
`define LDA_DP		12'h096
`define STA_DP		12'h097
`define EORA_DP		12'h098
`define ADCA_DP		12'h099
`define ORA_DP		12'h09A
`define ADDA_DP		12'h09B
`define CMPX_DP		12'h09C
`define JSR_DP		12'h09D
`define LDX_DP		12'h09E
`define STX_DP		12'h09F

`define SUBA_NDX	12'h0A0
`define CMPA_NDX	12'h0A1
`define SBCA_NDX	12'h0A2
`define SUBD_NDX	12'h0A3
`define ANDA_NDX	12'h0A4
`define BITA_NDX	12'h0A5
`define LDA_NDX		12'h0A6
`define STA_NDX		12'h0A7
`define EORA_NDX	12'h0A8
`define ADCA_NDX	12'h0A9
`define ORA_NDX		12'h0AA
`define ADDA_NDX	12'h0AB
`define CMPX_NDX	12'h0AC
`define JSR_NDX		12'h0AD
`define LDX_NDX		12'h0AE
`define STX_NDX		12'h0AF

`define SUBA_EXT	12'h0B0
`define CMPA_EXT	12'h0B1
`define SBCA_EXT	12'h0B2
`define SUBD_EXT	12'h0B3
`define ANDA_EXT	12'h0B4
`define BITA_EXT	12'h0B5
`define LDA_EXT		12'h0B6
`define STA_EXT		12'h0B7
`define EORA_EXT	12'h0B8
`define ADCA_EXT	12'h0B9
`define ORA_EXT		12'h0BA
`define ADDA_EXT	12'h0BB
`define CMPX_EXT	12'h0BC
`define JSR_EXT		12'h0BD
`define LDX_EXT		12'h0BE
`define STX_EXT		12'h0BF

`define SUBB_IMM	12'h0C0
`define CMPB_IMM	12'h0C1
`define SBCB_IMM	12'h0C2
`define ADDD_IMM	12'h0C3
`define ANDB_IMM	12'h0C4
`define BITB_IMM	12'h0C5
`define LDB_IMM		12'h0C6
`define EORB_IMM	12'h0C8
`define ADCB_IMM	12'h0C9
`define ORB_IMM		12'h0CA
`define ADDB_IMM	12'h0CB
`define LDD_IMM		12'h0CC
`define LDQ_IMM		12'h0CD
`define LDU_IMM		12'h0CE
`define JSR_FAR		12'h0CF

`define SUBB_DP		12'h0D0
`define CMPB_DP		12'h0D1
`define SBCB_DP		12'h0D2
`define ADDD_DP		12'h0D3
`define ANDB_DP		12'h0D4
`define BITB_DP		12'h0D5
`define LDB_DP		12'h0D6
`define STB_DP		12'h0D7
`define EORB_DP		12'h0D8
`define ADCB_DP		12'h0D9
`define ORB_DP		12'h0DA
`define ADDB_DP		12'h0DB
`define LDD_DP		12'h0DC
`define STD_DP		12'h0DD
`define LDU_DP		12'h0DE
`define STU_DP		12'h0DF

`define SUBB_NDX	12'h0E0
`define CMPB_NDX	12'h0E1
`define SBCB_NDX	12'h0E2
`define ADDD_NDX	12'h0E3
`define ANDB_NDX	12'h0E4
`define BITB_NDX	12'h0E5
`define LDB_NDX		12'h0E6
`define STB_NDX		12'h0E7
`define EORB_NDX	12'h0E8
`define ADCB_NDX	12'h0E9
`define ORB_NDX		12'h0EA
`define ADDB_NDX	12'h0EB
`define LDD_NDX		12'h0EC
`define STD_NDX		12'h0ED
`define LDU_NDX		12'h0EE
`define STU_NDX		12'h0EF

`define SUBB_EXT	12'h0F0
`define CMPB_EXT	12'h0F1
`define SBCB_EXT	12'h0F2
`define ADDD_EXT	12'h0F3
`define ANDB_EXT	12'h0F4
`define BITB_EXT	12'h0F5
`define LDB_EXT		12'h0F6
`define STB_EXT		12'h0F7
`define EORB_EXT	12'h0F8
`define ADCB_EXT	12'h0F9
`define ORB_EXT		12'h0FA
`define ADDB_EXT	12'h0FB
`define LDD_EXT		12'h0FC
`define STD_EXT		12'h0FD
`define LDU_EXT		12'h0FE
`define STU_EXT		12'h0FF

`define TFS			12'h11E
`define TTS			12'h11F

`define LBRN		12'h121
`define LBHI		12'h122
`define LBLS		12'h123
`define LBHS		12'h124
`define LBLO		12'h125
`define LBNE		12'h126
`define LBEQ		12'h127
`define LBVC		12'h128
`define LBVS		12'h129
`define LBPL		12'h12A
`define LBMI		12'h12B
`define LBGE		12'h12C
`define LBLT		12'h12D
`define LBGT		12'h12E
`define LBLE		12'h12F

`define SWI2		12'h13F
`define ASLD		12'h148
`define TSTD		12'h14D
`define SBCD_IMM	12'h182
`define CMPD_IMM	12'h183
`define ANDD_IMM	12'h184
`define ADCD_IMM	12'h189
`define CMPY_IMM	12'h18C
`define LDY_IMM		12'h18E
`define SBCD_DP		12'h192
`define CMPD_DP		12'h193
`define ANDD_DP		12'h194
`define ADCD_DP		12'h199
`define CMPY_DP		12'h19C
`define LDY_DP		12'h19E
`define STY_DP		12'h19F
`define SBCD_NDX	12'h1A2
`define CMPD_NDX	12'h1A3
`define ANDD_NDX	12'h1A4
`define ADCD_NDX	12'h1A9
`define CMPY_NDX	12'h1AC
`define LDY_NDX		12'h1AE
`define STY_NDX		12'h1AF
`define SBCD_EXT	12'h1B2
`define CMPD_EXT	12'h1B3
`define ANDD_EXT	12'h1B4
`define ADCD_EXT	12'h1B9
`define CMPY_EXT	12'h1BC
`define LDY_EXT		12'h1BE
`define STY_EXT		12'h1BF
`define LDS_IMM		12'h1CE
`define LDQ_DP		12'h1DC
`define STQ_DP		12'h1DD
`define LDS_DP		12'h1DE
`define STS_DP		12'h1DF
`define LDQ_NDX		12'h1EC
`define STQ_NDX		12'h1ED
`define LDS_NDX		12'h1EE
`define STS_NDX		12'h1EF
`define LDQ_EXT		12'h1FC
`define STQ_EXT		12'h1FD
`define LDS_EXT		12'h1FE
`define STS_EXT		12'h1FF
`define LDMD		12'h23D
`define SWI3		12'h23F
`define CMPU_IMM	12'h283
`define CMPS_IMM	12'h28C
`define CMPU_DP		12'h293
`define CMPS_DP		12'h29C
`define CMPU_NDX	12'h2A3
`define CMPS_NDX	12'h2AC
`define CMPU_EXT	12'h2B3
`define CMPS_EXT	12'h2BC

// Unused opcode
`define INT			12'h33E

`define LW_CCR		6'd0
`define LW_ACCA		6'd1
`define LW_ACCB		6'd2
`define LW_DPR		6'd3
`define LW_XH		6'd4
`define LW_XL		6'd5
`define LW_YH		6'd6
`define LW_YL		6'd7
`define LW_USPH		6'd8
`define LW_USPL		6'd9
`define LW_SSPH		6'd10
`define LW_SSPL		6'd11
`define LW_PCH		6'd12
`define LW_PCL		6'd13
`define LW_BL		6'd14
`define LW_BH		6'd15
`define LW_IAL		6'd16
`define LW_IAH		6'd17
`define LW_PC3124	6'd18
`define LW_PC2316	6'd19
`define LW_IA3124	6'd20
`define LW_IA2316	6'd21
`define LW_B3124	6'd22
`define LW_B2316	6'd23
`define LW_X3124	6'd24
`define LW_X2316	6'd25
`define LW_Y3124	6'd26
`define LW_Y2316	6'd27
`define LW_USP3124	6'd28
`define LW_USP2316	6'd29
`define LW_SSP3124	6'd30
`define LW_SSP2316	6'd31
`define LW_NOTHING	6'd63

`define SW_ACCDH	6'd0
`define SW_ACCDL	6'd1
`define SW_ACCA		6'd2
`define SW_ACCB		6'd3
`define SW_DPR		6'd4
`define SW_XL		6'd5
`define SW_XH		6'd6
`define SW_YL		6'd7
`define SW_YH		6'd8
`define SW_USPL		6'd9
`define SW_USPH		6'd10
`define SW_SSPL		6'd11
`define SW_SSPH		6'd12
`define SW_PCH		6'd13
`define SW_PCL		6'd14
`define SW_CCR		6'd15
`define SW_RES8		6'd16
`define SW_RES16L	6'd17
`define SW_RES16H	6'd18
`define SW_DEF8		6'd19
`define SW_PC3124	6'd20
`define SW_PC2316	6'd21
`define SW_ACCQ3124	6'd22
`define SW_ACCQ2316	6'd23
`define SW_ACCQ158	6'd24
`define SW_ACCQ70	6'd25
`define SW_X3124	6'd26
`define SW_X2316	6'd27
`define SW_Y3124	6'd28
`define SW_Y2316	6'd29
`define SW_USP3124	6'd30
`define SW_USP2316	6'd31
`define SW_SSP3124	6'd32
`define SW_SSP2316	6'd33
`define SW_ACCA3124 6'd34
`define SW_ACCA2316 6'd35
`define SW_ACCA158 	6'd36
`define SW_ACCA70	6'd37
`define SW_ACCB3124 6'd38
`define SW_ACCB2316 6'd39
`define SW_ACCB158 	6'd40
`define SW_ACCB70	6'd41
`define SW_NOTHING	6'd63

endpackage
