
module 