package const_pkg;

`define TRUE	1
`define FALSE	0
`define HIGH	1
`define LOW		0
`define VAL		1
`define INV		0

 parameter TRUE = `TRUE;
 parameter FALSE = `FALSE;
 parameter VAL = `VAL;
 parameter INV = `INV;
 parameter HIGH = `HIGH;
 parameter LOW = `LOW;

endpackage
