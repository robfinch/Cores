rommem[0] <= 16'hFF40;
rommem[1] <= 16'h1000;
rommem[2] <= 16'hFFFC;
rommem[3] <= 16'h0010;
rommem[4] <= 16'h4141;
rommem[5] <= 16'h3030;
rommem[6] <= 16'h3030;
rommem[7] <= 16'h3030;
rommem[8] <= 16'h33FC;
rommem[9] <= 16'hA1A1;
rommem[10] <= 16'hFFDC;
rommem[11] <= 16'h0600;
rommem[12] <= 16'h7000;
rommem[13] <= 16'h7200;
rommem[14] <= 16'h7400;
rommem[15] <= 16'h7600;
rommem[16] <= 16'h7800;
rommem[17] <= 16'h7A00;
rommem[18] <= 16'h7C00;
rommem[19] <= 16'h7E00;
rommem[20] <= 16'h4288;
rommem[21] <= 16'h4289;
rommem[22] <= 16'h428A;
rommem[23] <= 16'h428B;
rommem[24] <= 16'h428C;
rommem[25] <= 16'h428D;
rommem[26] <= 16'h428E;
rommem[27] <= 16'h4E67;
rommem[28] <= 16'h6100;
rommem[29] <= 16'h134E;
rommem[30] <= 16'h33FC;
rommem[31] <= 16'hA2A2;
rommem[32] <= 16'hFFDC;
rommem[33] <= 16'h0600;
rommem[34] <= 16'h13FC;
rommem[35] <= 16'h0028;
rommem[36] <= 16'h0001;
rommem[37] <= 16'h041B;
rommem[38] <= 16'h13FC;
rommem[39] <= 16'h0020;
rommem[40] <= 16'h0001;
rommem[41] <= 16'h041A;
rommem[42] <= 16'h4239;
rommem[43] <= 16'h0001;
rommem[44] <= 16'h0419;
rommem[45] <= 16'h4239;
rommem[46] <= 16'h0001;
rommem[47] <= 16'h0418;
rommem[48] <= 16'h4279;
rommem[49] <= 16'h0001;
rommem[50] <= 16'h041C;
rommem[51] <= 16'h23FC;
rommem[52] <= 16'h0002;
rommem[53] <= 16'h0000;
rommem[54] <= 16'h0001;
rommem[55] <= 16'h0420;
rommem[56] <= 16'h6100;
rommem[57] <= 16'h03E8;
rommem[58] <= 16'h6100;
rommem[59] <= 16'h03FC;
rommem[60] <= 16'h4DF9;
rommem[61] <= 16'hFFDC;
rommem[62] <= 16'h0000;
rommem[63] <= 16'h426E;
rommem[64] <= 16'h0C06;
rommem[65] <= 16'h2D7C;
rommem[66] <= 16'h8888;
rommem[67] <= 16'h8888;
rommem[68] <= 16'h0C08;
rommem[69] <= 16'h2D7C;
rommem[70] <= 16'h0123;
rommem[71] <= 16'h4567;
rommem[72] <= 16'h0C0C;
rommem[73] <= 16'h6100;
rommem[74] <= 16'h02BC;
rommem[75] <= 16'h33FC;
rommem[76] <= 16'hA2A2;
rommem[77] <= 16'hFFDC;
rommem[78] <= 16'h0600;
rommem[79] <= 16'h2A7C;
rommem[80] <= 16'hFFE0;
rommem[81] <= 16'h0000;
rommem[82] <= 16'h3B7C;
rommem[83] <= 16'h4000;
rommem[84] <= 16'h0584;
rommem[85] <= 16'h6100;
rommem[86] <= 16'h1186;
rommem[87] <= 16'h6100;
rommem[88] <= 16'h1222;
rommem[89] <= 16'h6100;
rommem[90] <= 16'h02B2;
rommem[91] <= 16'h33FC;
rommem[92] <= 16'hA3A3;
rommem[93] <= 16'hFFDC;
rommem[94] <= 16'h0600;
rommem[95] <= 16'h33FC;
rommem[96] <= 16'h7FFF;
rommem[97] <= 16'h0001;
rommem[98] <= 16'h0002;
rommem[99] <= 16'h33FC;
rommem[100] <= 16'h000F;
rommem[101] <= 16'h0001;
rommem[102] <= 16'h0004;
rommem[103] <= 16'h41F9;
rommem[104] <= 16'hFFFC;
rommem[105] <= 16'h168B;
rommem[106] <= 16'h7200;
rommem[107] <= 16'h7400;
rommem[108] <= 16'h6100;
rommem[109] <= 16'h03D6;
rommem[110] <= 16'h33FC;
rommem[111] <= 16'hA4A4;
rommem[112] <= 16'hFFDC;
rommem[113] <= 16'h0600;
rommem[114] <= 16'h47F9;
rommem[115] <= 16'hFFFC;
rommem[116] <= 16'h00EE;
rommem[117] <= 16'h6000;
rommem[118] <= 16'h0FD8;
rommem[119] <= 16'h60FE;
rommem[120] <= 16'h2F01;
rommem[121] <= 16'h123C;
rommem[122] <= 16'h000D;
rommem[123] <= 16'h4EB9;
rommem[124] <= 16'hFFFC;
rommem[125] <= 16'h013A;
rommem[126] <= 16'h123C;
rommem[127] <= 16'h000A;
rommem[128] <= 16'h4EB9;
rommem[129] <= 16'hFFFC;
rommem[130] <= 16'h013A;
rommem[131] <= 16'h221F;
rommem[132] <= 16'h4E75;
rommem[133] <= 16'h1039;
rommem[134] <= 16'h0001;
rommem[135] <= 16'h0418;
rommem[136] <= 16'h0240;
rommem[137] <= 16'h007F;
rommem[138] <= 16'h1439;
rommem[139] <= 16'h0001;
rommem[140] <= 16'h041B;
rommem[141] <= 16'h4882;
rommem[142] <= 16'hC0C2;
rommem[143] <= 16'h1439;
rommem[144] <= 16'h0001;
rommem[145] <= 16'h0419;
rommem[146] <= 16'h0242;
rommem[147] <= 16'h00FF;
rommem[148] <= 16'hD042;
rommem[149] <= 16'h33C0;
rommem[150] <= 16'h0001;
rommem[151] <= 16'h041C;
rommem[152] <= 16'hD0B9;
rommem[153] <= 16'h0001;
rommem[154] <= 16'h0420;
rommem[155] <= 16'h2040;
rommem[156] <= 16'h4E75;
rommem[157] <= 16'h0C01;
rommem[158] <= 16'h000D;
rommem[159] <= 16'h6608;
rommem[160] <= 16'h4239;
rommem[161] <= 16'h0001;
rommem[162] <= 16'h0419;
rommem[163] <= 16'h4E75;
rommem[164] <= 16'h0C01;
rommem[165] <= 16'h0091;
rommem[166] <= 16'h6616;
rommem[167] <= 16'h0C39;
rommem[168] <= 16'h004F;
rommem[169] <= 16'h0001;
rommem[170] <= 16'h0419;
rommem[171] <= 16'h670A;
rommem[172] <= 16'h5239;
rommem[173] <= 16'h0001;
rommem[174] <= 16'h0419;
rommem[175] <= 16'h6000;
rommem[176] <= 16'h02C4;
rommem[177] <= 16'h4E75;
rommem[178] <= 16'h0C01;
rommem[179] <= 16'h0090;
rommem[180] <= 16'h6614;
rommem[181] <= 16'h0C39;
rommem[182] <= 16'h0000;
rommem[183] <= 16'h0001;
rommem[184] <= 16'h0418;
rommem[185] <= 16'h67EE;
rommem[186] <= 16'h5339;
rommem[187] <= 16'h0001;
rommem[188] <= 16'h0418;
rommem[189] <= 16'h6000;
rommem[190] <= 16'h02A8;
rommem[191] <= 16'h0C01;
rommem[192] <= 16'h0093;
rommem[193] <= 16'h6614;
rommem[194] <= 16'h0C39;
rommem[195] <= 16'h0000;
rommem[196] <= 16'h0001;
rommem[197] <= 16'h0419;
rommem[198] <= 16'h67D4;
rommem[199] <= 16'h5339;
rommem[200] <= 16'h0001;
rommem[201] <= 16'h0419;
rommem[202] <= 16'h6000;
rommem[203] <= 16'h028E;
rommem[204] <= 16'h0C01;
rommem[205] <= 16'h0092;
rommem[206] <= 16'h6614;
rommem[207] <= 16'h0C39;
rommem[208] <= 16'h003F;
rommem[209] <= 16'h0001;
rommem[210] <= 16'h0418;
rommem[211] <= 16'h67BA;
rommem[212] <= 16'h5279;
rommem[213] <= 16'h0001;
rommem[214] <= 16'h0418;
rommem[215] <= 16'h6000;
rommem[216] <= 16'h0274;
rommem[217] <= 16'h0C01;
rommem[218] <= 16'h0094;
rommem[219] <= 16'h661E;
rommem[220] <= 16'h0C39;
rommem[221] <= 16'h0000;
rommem[222] <= 16'h0001;
rommem[223] <= 16'h0419;
rommem[224] <= 16'h670A;
rommem[225] <= 16'h4239;
rommem[226] <= 16'h0001;
rommem[227] <= 16'h0419;
rommem[228] <= 16'h6000;
rommem[229] <= 16'h025A;
rommem[230] <= 16'h4239;
rommem[231] <= 16'h0001;
rommem[232] <= 16'h0418;
rommem[233] <= 16'h6000;
rommem[234] <= 16'h0250;
rommem[235] <= 16'h48E7;
rommem[236] <= 16'hE080;
rommem[237] <= 16'h0C01;
rommem[238] <= 16'h0099;
rommem[239] <= 16'h660C;
rommem[240] <= 16'h6100;
rommem[241] <= 16'hFF28;
rommem[242] <= 16'h1039;
rommem[243] <= 16'h0001;
rommem[244] <= 16'h0419;
rommem[245] <= 16'h6020;
rommem[246] <= 16'h0C01;
rommem[247] <= 16'h0000;
rommem[248] <= 16'h6632;
rommem[249] <= 16'h0C39;
rommem[250] <= 16'h0000;
rommem[251] <= 16'h0001;
rommem[252] <= 16'h0419;
rommem[253] <= 16'h6752;
rommem[254] <= 16'h5339;
rommem[255] <= 16'h0001;
rommem[256] <= 16'h0419;
rommem[257] <= 16'h6100;
rommem[258] <= 16'hFF06;
rommem[259] <= 16'h1039;
rommem[260] <= 16'h0001;
rommem[261] <= 16'h0419;
rommem[262] <= 16'h10E8;
rommem[263] <= 16'h0001;
rommem[264] <= 16'h5200;
rommem[265] <= 16'hB039;
rommem[266] <= 16'h0001;
rommem[267] <= 16'h041B;
rommem[268] <= 16'h65F2;
rommem[269] <= 16'h103C;
rommem[270] <= 16'h0020;
rommem[271] <= 16'h1140;
rommem[272] <= 16'hFFFF;
rommem[273] <= 16'h602A;
rommem[274] <= 16'h0C01;
rommem[275] <= 16'h000A;
rommem[276] <= 16'h671C;
rommem[277] <= 16'h6100;
rommem[278] <= 16'hFEDE;
rommem[279] <= 16'h1081;
rommem[280] <= 16'h1001;
rommem[281] <= 16'h4880;
rommem[282] <= 16'h6100;
rommem[283] <= 16'h0194;
rommem[284] <= 16'h6100;
rommem[285] <= 16'h001A;
rommem[286] <= 16'h6100;
rommem[287] <= 16'h01E6;
rommem[288] <= 16'h4CDF;
rommem[289] <= 16'h0107;
rommem[290] <= 16'h4E75;
rommem[291] <= 16'h6100;
rommem[292] <= 16'h002C;
rommem[293] <= 16'h6100;
rommem[294] <= 16'h01D8;
rommem[295] <= 16'h4CDF;
rommem[296] <= 16'h0107;
rommem[297] <= 16'h4E75;
rommem[298] <= 16'h5279;
rommem[299] <= 16'h0001;
rommem[300] <= 16'h041C;
rommem[301] <= 16'h5239;
rommem[302] <= 16'h0001;
rommem[303] <= 16'h0419;
rommem[304] <= 16'h1039;
rommem[305] <= 16'h0001;
rommem[306] <= 16'h041B;
rommem[307] <= 16'hB039;
rommem[308] <= 16'h0001;
rommem[309] <= 16'h0419;
rommem[310] <= 16'h643A;
rommem[311] <= 16'h4239;
rommem[312] <= 16'h0001;
rommem[313] <= 16'h0419;
rommem[314] <= 16'h5239;
rommem[315] <= 16'h0001;
rommem[316] <= 16'h0418;
rommem[317] <= 16'h1039;
rommem[318] <= 16'h0001;
rommem[319] <= 16'h041A;
rommem[320] <= 16'hB039;
rommem[321] <= 16'h0001;
rommem[322] <= 16'h0418;
rommem[323] <= 16'h6220;
rommem[324] <= 16'h1039;
rommem[325] <= 16'h0001;
rommem[326] <= 16'h041A;
rommem[327] <= 16'h13C0;
rommem[328] <= 16'h0001;
rommem[329] <= 16'h0418;
rommem[330] <= 16'h5339;
rommem[331] <= 16'h0001;
rommem[332] <= 16'h0418;
rommem[333] <= 16'h4880;
rommem[334] <= 16'hE340;
rommem[335] <= 16'h9179;
rommem[336] <= 16'h0001;
rommem[337] <= 16'h041C;
rommem[338] <= 16'h6100;
rommem[339] <= 16'h0B76;
rommem[340] <= 16'h4E75;
rommem[341] <= 16'h48E7;
rommem[342] <= 16'hC040;
rommem[343] <= 16'h4281;
rommem[344] <= 16'h1219;
rommem[345] <= 16'h0C01;
rommem[346] <= 16'h0000;
rommem[347] <= 16'h6706;
rommem[348] <= 16'h6100;
rommem[349] <= 16'hFE80;
rommem[350] <= 16'h60F0;
rommem[351] <= 16'h4CDF;
rommem[352] <= 16'h0203;
rommem[353] <= 16'h4E75;
rommem[354] <= 16'h6100;
rommem[355] <= 16'hFFE4;
rommem[356] <= 16'h6000;
rommem[357] <= 16'hFE26;
rommem[358] <= 16'h48E7;
rommem[359] <= 16'hC040;
rommem[360] <= 16'h0241;
rommem[361] <= 16'h00FF;
rommem[362] <= 16'h2001;
rommem[363] <= 16'h1219;
rommem[364] <= 16'h0C01;
rommem[365] <= 16'h0000;
rommem[366] <= 16'h6708;
rommem[367] <= 16'h6100;
rommem[368] <= 16'hFE5A;
rommem[369] <= 16'h57C8;
rommem[370] <= 16'hFFF2;
rommem[371] <= 16'h4CDF;
rommem[372] <= 16'h0203;
rommem[373] <= 16'h4E75;
rommem[374] <= 16'h6100;
rommem[375] <= 16'hFFDE;
rommem[376] <= 16'h6000;
rommem[377] <= 16'hFDFE;
rommem[378] <= 16'h0C41;
rommem[379] <= 16'h00FF;
rommem[380] <= 16'h670E;
rommem[381] <= 16'h0C41;
rommem[382] <= 16'hFF00;
rommem[383] <= 16'h6718;
rommem[384] <= 16'h4EB9;
rommem[385] <= 16'hFFFC;
rommem[386] <= 16'h0DDC;
rommem[387] <= 16'h4E75;
rommem[388] <= 16'h1239;
rommem[389] <= 16'h0001;
rommem[390] <= 16'h0419;
rommem[391] <= 16'hE141;
rommem[392] <= 16'h1239;
rommem[393] <= 16'h0001;
rommem[394] <= 16'h0418;
rommem[395] <= 16'h4E75;
rommem[396] <= 16'h48E7;
rommem[397] <= 16'h6000;
rommem[398] <= 16'h13C1;
rommem[399] <= 16'h0001;
rommem[400] <= 16'h0418;
rommem[401] <= 16'hE049;
rommem[402] <= 16'h13C1;
rommem[403] <= 16'h0001;
rommem[404] <= 16'h0419;
rommem[405] <= 16'h1239;
rommem[406] <= 16'h0001;
rommem[407] <= 16'h0418;
rommem[408] <= 16'h4881;
rommem[409] <= 16'h1439;
rommem[410] <= 16'h0001;
rommem[411] <= 16'h041B;
rommem[412] <= 16'h4882;
rommem[413] <= 16'hC2C2;
rommem[414] <= 16'h1439;
rommem[415] <= 16'h0001;
rommem[416] <= 16'h0419;
rommem[417] <= 16'hD242;
rommem[418] <= 16'h33C1;
rommem[419] <= 16'h0001;
rommem[420] <= 16'h041C;
rommem[421] <= 16'h4CDF;
rommem[422] <= 16'h0006;
rommem[423] <= 16'h4E75;
rommem[424] <= 16'h207C;
rommem[425] <= 16'hFF80;
rommem[426] <= 16'h0000;
rommem[427] <= 16'h700F;
rommem[428] <= 16'h223C;
rommem[429] <= 16'h0001;
rommem[430] <= 16'h4000;
rommem[431] <= 16'h30C0;
rommem[432] <= 16'h5381;
rommem[433] <= 16'h66FA;
rommem[434] <= 16'h4E75;
rommem[435] <= 16'h33FC;
rommem[436] <= 16'h0707;
rommem[437] <= 16'h0001;
rommem[438] <= 16'h0006;
rommem[439] <= 16'h41F9;
rommem[440] <= 16'hFFFC;
rommem[441] <= 16'h16A3;
rommem[442] <= 16'h223C;
rommem[443] <= 16'h0000;
rommem[444] <= 16'h1000;
rommem[445] <= 16'h227C;
rommem[446] <= 16'hFF8B;
rommem[447] <= 16'h8000;
rommem[448] <= 16'h7000;
rommem[449] <= 16'h1018;
rommem[450] <= 16'h32C0;
rommem[451] <= 16'h51C9;
rommem[452] <= 16'hFFFA;
rommem[453] <= 16'h4E75;
rommem[454] <= 16'h2C7C;
rommem[455] <= 16'hFFE0;
rommem[456] <= 16'h0000;
rommem[457] <= 16'h4840;
rommem[458] <= 16'h302E;
rommem[459] <= 16'h042C;
rommem[460] <= 16'hB07C;
rommem[461] <= 16'h001C;
rommem[462] <= 16'h64F6;
rommem[463] <= 16'h4840;
rommem[464] <= 16'h3D40;
rommem[465] <= 16'h0420;
rommem[466] <= 16'h3D79;
rommem[467] <= 16'h0001;
rommem[468] <= 16'h0002;
rommem[469] <= 16'h0422;
rommem[470] <= 16'h3D79;
rommem[471] <= 16'h0001;
rommem[472] <= 16'h0004;
rommem[473] <= 16'h0424;
rommem[474] <= 16'h3D41;
rommem[475] <= 16'h0426;
rommem[476] <= 16'h3D42;
rommem[477] <= 16'h0428;
rommem[478] <= 16'h3D7C;
rommem[479] <= 16'h0707;
rommem[480] <= 16'h042A;
rommem[481] <= 16'h3D7C;
rommem[482] <= 16'h0000;
rommem[483] <= 16'h042E;
rommem[484] <= 16'h4E75;
rommem[485] <= 16'h48E7;
rommem[486] <= 16'h4002;
rommem[487] <= 16'h2C7C;
rommem[488] <= 16'hFFE0;
rommem[489] <= 16'h0000;
rommem[490] <= 16'h4840;
rommem[491] <= 16'h302E;
rommem[492] <= 16'h042C;
rommem[493] <= 16'hB07C;
rommem[494] <= 16'h001C;
rommem[495] <= 16'h64F6;
rommem[496] <= 16'h4840;
rommem[497] <= 16'h3D40;
rommem[498] <= 16'h0420;
rommem[499] <= 16'h3D79;
rommem[500] <= 16'h0001;
rommem[501] <= 16'h0002;
rommem[502] <= 16'h0422;
rommem[503] <= 16'h3D79;
rommem[504] <= 16'h0001;
rommem[505] <= 16'h0004;
rommem[506] <= 16'h0424;
rommem[507] <= 16'h1239;
rommem[508] <= 16'h0001;
rommem[509] <= 16'h0419;
rommem[510] <= 16'h4881;
rommem[511] <= 16'hE741;
rommem[512] <= 16'h3D41;
rommem[513] <= 16'h0426;
rommem[514] <= 16'h1239;
rommem[515] <= 16'h0001;
rommem[516] <= 16'h0418;
rommem[517] <= 16'h4881;
rommem[518] <= 16'hE741;
rommem[519] <= 16'h3D41;
rommem[520] <= 16'h0428;
rommem[521] <= 16'h3D7C;
rommem[522] <= 16'h0707;
rommem[523] <= 16'h042A;
rommem[524] <= 16'h3D7C;
rommem[525] <= 16'h0000;
rommem[526] <= 16'h042E;
rommem[527] <= 16'h4CDF;
rommem[528] <= 16'h4002;
rommem[529] <= 16'h4E75;
rommem[530] <= 16'h48E7;
rommem[531] <= 16'h4002;
rommem[532] <= 16'h2C7C;
rommem[533] <= 16'hFFE0;
rommem[534] <= 16'h0000;
rommem[535] <= 16'h3D7C;
rommem[536] <= 16'h0A0A;
rommem[537] <= 16'h0444;
rommem[538] <= 16'h1239;
rommem[539] <= 16'h0001;
rommem[540] <= 16'h0419;
rommem[541] <= 16'h4881;
rommem[542] <= 16'hE741;
rommem[543] <= 16'h5341;
rommem[544] <= 16'h3D41;
rommem[545] <= 16'h0440;
rommem[546] <= 16'h1239;
rommem[547] <= 16'h0001;
rommem[548] <= 16'h0418;
rommem[549] <= 16'h4881;
rommem[550] <= 16'hE741;
rommem[551] <= 16'h5341;
rommem[552] <= 16'h3D41;
rommem[553] <= 16'h0442;
rommem[554] <= 16'h4CDF;
rommem[555] <= 16'h4002;
rommem[556] <= 16'h4E75;
rommem[557] <= 16'h2F0E;
rommem[558] <= 16'h2C7C;
rommem[559] <= 16'hFFE0;
rommem[560] <= 16'h0000;
rommem[561] <= 16'h3D7C;
rommem[562] <= 16'h7FFF;
rommem[563] <= 16'h0446;
rommem[564] <= 16'h3D7C;
rommem[565] <= 16'h0004;
rommem[566] <= 16'h0448;
rommem[567] <= 16'h2C5F;
rommem[568] <= 16'h4E75;
rommem[569] <= 16'h48E7;
rommem[570] <= 16'h4082;
rommem[571] <= 16'h41F9;
rommem[572] <= 16'hFFFC;
rommem[573] <= 16'h0490;
rommem[574] <= 16'h2C7C;
rommem[575] <= 16'hFFE0;
rommem[576] <= 16'h0460;
rommem[577] <= 16'h720F;
rommem[578] <= 16'h3CD8;
rommem[579] <= 16'h51C9;
rommem[580] <= 16'hFFFC;
rommem[581] <= 16'h4CDF;
rommem[582] <= 16'h4102;
rommem[583] <= 16'h4E75;
rommem[584] <= 16'h03FF;
rommem[585] <= 16'h0201;
rommem[586] <= 16'h0201;
rommem[587] <= 16'h0201;
rommem[588] <= 16'h0201;
rommem[589] <= 16'h0201;
rommem[590] <= 16'h0201;
rommem[591] <= 16'h0201;
rommem[592] <= 16'h0231;
rommem[593] <= 16'h03FF;
rommem[594] <= 16'h0000;
rommem[595] <= 16'h0000;
rommem[596] <= 16'h0000;
rommem[597] <= 16'h0000;
rommem[598] <= 16'h0000;
rommem[599] <= 16'h0000;
rommem[600] <= 16'h7000;
rommem[601] <= 16'h1018;
rommem[602] <= 16'h6708;
rommem[603] <= 16'h6100;
rommem[604] <= 16'hFED4;
rommem[605] <= 16'h5041;
rommem[606] <= 16'h60F2;
rommem[607] <= 16'h4E75;
rommem[608] <= 16'h3F01;
rommem[609] <= 16'h0201;
rommem[610] <= 16'h000F;
rommem[611] <= 16'h0601;
rommem[612] <= 16'h0030;
rommem[613] <= 16'h0C01;
rommem[614] <= 16'h0039;
rommem[615] <= 16'h6302;
rommem[616] <= 16'h5E01;
rommem[617] <= 16'h6100;
rommem[618] <= 16'hFC66;
rommem[619] <= 16'h321F;
rommem[620] <= 16'h4E75;
rommem[621] <= 16'h3F01;
rommem[622] <= 16'hE819;
rommem[623] <= 16'h6100;
rommem[624] <= 16'hFFE0;
rommem[625] <= 16'hE919;
rommem[626] <= 16'h6100;
rommem[627] <= 16'hFFDA;
rommem[628] <= 16'h321F;
rommem[629] <= 16'h4E75;
rommem[630] <= 16'hE199;
rommem[631] <= 16'h6100;
rommem[632] <= 16'hFFEA;
rommem[633] <= 16'hE199;
rommem[634] <= 16'h6100;
rommem[635] <= 16'hFFE4;
rommem[636] <= 16'hE199;
rommem[637] <= 16'h6100;
rommem[638] <= 16'hFFDE;
rommem[639] <= 16'hE199;
rommem[640] <= 16'h6100;
rommem[641] <= 16'hFFD8;
rommem[642] <= 16'h4E75;
rommem[643] <= 16'h123C;
rommem[644] <= 16'h003A;
rommem[645] <= 16'h4EB9;
rommem[646] <= 16'hFFFC;
rommem[647] <= 16'h013A;
rommem[648] <= 16'h2208;
rommem[649] <= 16'h4EB9;
rommem[650] <= 16'hFFFC;
rommem[651] <= 16'h04EC;
rommem[652] <= 16'h7407;
rommem[653] <= 16'h123C;
rommem[654] <= 16'h0020;
rommem[655] <= 16'h4EB9;
rommem[656] <= 16'hFFFC;
rommem[657] <= 16'h013A;
rommem[658] <= 16'h1218;
rommem[659] <= 16'h4EB9;
rommem[660] <= 16'hFFFC;
rommem[661] <= 16'h04DA;
rommem[662] <= 16'h51CA;
rommem[663] <= 16'hFFEC;
rommem[664] <= 16'h4EF9;
rommem[665] <= 16'hFFFC;
rommem[666] <= 16'h00F0;
rommem[667] <= 16'h1239;
rommem[668] <= 16'hFFDC;
rommem[669] <= 16'h0001;
rommem[670] <= 16'h4E75;
rommem[671] <= 16'h7200;
rommem[672] <= 16'h1239;
rommem[673] <= 16'hFFDC;
rommem[674] <= 16'h0000;
rommem[675] <= 16'h13FC;
rommem[676] <= 16'h0000;
rommem[677] <= 16'hFFDC;
rommem[678] <= 16'h0001;
rommem[679] <= 16'h4E75;
rommem[680] <= 16'h2F03;
rommem[681] <= 16'h363C;
rommem[682] <= 16'h0064;
rommem[683] <= 16'h6100;
rommem[684] <= 16'hFFDE;
rommem[685] <= 16'h4A01;
rommem[686] <= 16'h6B0E;
rommem[687] <= 16'h6100;
rommem[688] <= 16'h02C4;
rommem[689] <= 16'h51CB;
rommem[690] <= 16'hFFF2;
rommem[691] <= 16'h261F;
rommem[692] <= 16'h72FF;
rommem[693] <= 16'h4E75;
rommem[694] <= 16'h6100;
rommem[695] <= 16'hFFD0;
rommem[696] <= 16'h261F;
rommem[697] <= 16'h4E75;
rommem[698] <= 16'h48E7;
rommem[699] <= 16'h3000;
rommem[700] <= 16'h7664;
rommem[701] <= 16'h6100;
rommem[702] <= 16'hFFBA;
rommem[703] <= 16'h0801;
rommem[704] <= 16'h0006;
rommem[705] <= 16'h6610;
rommem[706] <= 16'h6100;
rommem[707] <= 16'h029E;
rommem[708] <= 16'h51CB;
rommem[709] <= 16'hFFF0;
rommem[710] <= 16'h4CDF;
rommem[711] <= 16'h000C;
rommem[712] <= 16'h72FF;
rommem[713] <= 16'h4E75;
rommem[714] <= 16'h4CDF;
rommem[715] <= 16'h000C;
rommem[716] <= 16'h7200;
rommem[717] <= 16'h4E75;
rommem[718] <= 16'h1239;
rommem[719] <= 16'hFFDC;
rommem[720] <= 16'h0001;
rommem[721] <= 16'h6A06;
rommem[722] <= 16'h123C;
rommem[723] <= 16'h0001;
rommem[724] <= 16'h4E75;
rommem[725] <= 16'h4201;
rommem[726] <= 16'h4E75;
rommem[727] <= 16'h6100;
rommem[728] <= 16'h0022;
rommem[729] <= 16'h0C39;
rommem[730] <= 16'h0000;
rommem[731] <= 16'h0001;
rommem[732] <= 16'h0424;
rommem[733] <= 16'h670C;
rommem[734] <= 16'h0C01;
rommem[735] <= 16'h000D;
rommem[736] <= 16'h6700;
rommem[737] <= 16'hFB2E;
rommem[738] <= 16'h6100;
rommem[739] <= 16'hFB74;
rommem[740] <= 16'h4E75;
rommem[741] <= 16'h4239;
rommem[742] <= 16'h0001;
rommem[743] <= 16'h0425;
rommem[744] <= 16'h6008;
rommem[745] <= 16'h13FC;
rommem[746] <= 16'hFFFF;
rommem[747] <= 16'h0001;
rommem[748] <= 16'h0425;
rommem[749] <= 16'h48E7;
rommem[750] <= 16'h3080;
rommem[751] <= 16'h6100;
rommem[752] <= 16'hFF56;
rommem[753] <= 16'h6B10;
rommem[754] <= 16'h4A39;
rommem[755] <= 16'h0001;
rommem[756] <= 16'h0425;
rommem[757] <= 16'h6BF2;
rommem[758] <= 16'h4CDF;
rommem[759] <= 16'h010C;
rommem[760] <= 16'h72FF;
rommem[761] <= 16'h4E75;
rommem[762] <= 16'h6100;
rommem[763] <= 16'hFF48;
rommem[764] <= 16'h33FC;
rommem[765] <= 16'h0001;
rommem[766] <= 16'hFFDC;
rommem[767] <= 16'h0600;
rommem[768] <= 16'hB23C;
rommem[769] <= 16'h00F0;
rommem[770] <= 16'h6700;
rommem[771] <= 16'h00CA;
rommem[772] <= 16'hB23C;
rommem[773] <= 16'h00E0;
rommem[774] <= 16'h6700;
rommem[775] <= 16'h00CE;
rommem[776] <= 16'hB23C;
rommem[777] <= 16'h0014;
rommem[778] <= 16'h6700;
rommem[779] <= 16'h00D2;
rommem[780] <= 16'hB23C;
rommem[781] <= 16'h0012;
rommem[782] <= 16'h6700;
rommem[783] <= 16'h0134;
rommem[784] <= 16'hB23C;
rommem[785] <= 16'h0059;
rommem[786] <= 16'h6700;
rommem[787] <= 16'h012C;
rommem[788] <= 16'hB23C;
rommem[789] <= 16'h0077;
rommem[790] <= 16'h6700;
rommem[791] <= 16'h014C;
rommem[792] <= 16'hB23C;
rommem[793] <= 16'h0058;
rommem[794] <= 16'h6700;
rommem[795] <= 16'h0154;
rommem[796] <= 16'hB23C;
rommem[797] <= 16'h007E;
rommem[798] <= 16'h6700;
rommem[799] <= 16'h015C;
rommem[800] <= 16'hB23C;
rommem[801] <= 16'h0011;
rommem[802] <= 16'h6700;
rommem[803] <= 16'h00CA;
rommem[804] <= 16'h1439;
rommem[805] <= 16'h0001;
rommem[806] <= 16'h0426;
rommem[807] <= 16'h13FC;
rommem[808] <= 16'h0000;
rommem[809] <= 16'h0001;
rommem[810] <= 16'h0426;
rommem[811] <= 16'h4A02;
rommem[812] <= 16'h6684;
rommem[813] <= 16'hB23C;
rommem[814] <= 16'h000D;
rommem[815] <= 16'h6700;
rommem[816] <= 16'h00D8;
rommem[817] <= 16'h1439;
rommem[818] <= 16'h0001;
rommem[819] <= 16'h0427;
rommem[820] <= 16'h6A1E;
rommem[821] <= 16'h0202;
rommem[822] <= 16'h007F;
rommem[823] <= 16'h13C2;
rommem[824] <= 16'h0001;
rommem[825] <= 16'h0427;
rommem[826] <= 16'h13FC;
rommem[827] <= 16'h0000;
rommem[828] <= 16'h0001;
rommem[829] <= 16'h0426;
rommem[830] <= 16'h41F9;
rommem[831] <= 16'hFFFC;
rommem[832] <= 16'h0AB4;
rommem[833] <= 16'h1230;
rommem[834] <= 16'h1000;
rommem[835] <= 16'h603A;
rommem[836] <= 16'h0802;
rommem[837] <= 16'h0002;
rommem[838] <= 16'h6710;
rommem[839] <= 16'h0241;
rommem[840] <= 16'h007F;
rommem[841] <= 16'h41F9;
rommem[842] <= 16'hFFFC;
rommem[843] <= 16'h0A34;
rommem[844] <= 16'h1230;
rommem[845] <= 16'h1000;
rommem[846] <= 16'h6024;
rommem[847] <= 16'h0802;
rommem[848] <= 16'h0000;
rommem[849] <= 16'h670C;
rommem[850] <= 16'h41F9;
rommem[851] <= 16'hFFFC;
rommem[852] <= 16'h0934;
rommem[853] <= 16'h1230;
rommem[854] <= 16'h1000;
rommem[855] <= 16'h6012;
rommem[856] <= 16'h41F9;
rommem[857] <= 16'hFFFC;
rommem[858] <= 16'h0834;
rommem[859] <= 16'h1230;
rommem[860] <= 16'h1000;
rommem[861] <= 16'h33FC;
rommem[862] <= 16'h0202;
rommem[863] <= 16'hFFDC;
rommem[864] <= 16'h0600;
rommem[865] <= 16'h33FC;
rommem[866] <= 16'h0303;
rommem[867] <= 16'hFFDC;
rommem[868] <= 16'h0600;
rommem[869] <= 16'h4CDF;
rommem[870] <= 16'h010C;
rommem[871] <= 16'h4E75;
rommem[872] <= 16'h13FC;
rommem[873] <= 16'hFFFF;
rommem[874] <= 16'h0001;
rommem[875] <= 16'h0426;
rommem[876] <= 16'h6000;
rommem[877] <= 16'hFF04;
rommem[878] <= 16'h0039;
rommem[879] <= 16'h0080;
rommem[880] <= 16'h0001;
rommem[881] <= 16'h0427;
rommem[882] <= 16'h6000;
rommem[883] <= 16'hFEF8;
rommem[884] <= 16'h1239;
rommem[885] <= 16'h0001;
rommem[886] <= 16'h0426;
rommem[887] <= 16'h4239;
rommem[888] <= 16'h0001;
rommem[889] <= 16'h0426;
rommem[890] <= 16'h4A01;
rommem[891] <= 16'h6A0C;
rommem[892] <= 16'h08B9;
rommem[893] <= 16'h0002;
rommem[894] <= 16'h0001;
rommem[895] <= 16'h0427;
rommem[896] <= 16'h6000;
rommem[897] <= 16'hFEDC;
rommem[898] <= 16'h08F9;
rommem[899] <= 16'h0002;
rommem[900] <= 16'h0001;
rommem[901] <= 16'h0427;
rommem[902] <= 16'h6000;
rommem[903] <= 16'hFED0;
rommem[904] <= 16'h1239;
rommem[905] <= 16'h0001;
rommem[906] <= 16'h0426;
rommem[907] <= 16'h4239;
rommem[908] <= 16'h0001;
rommem[909] <= 16'h0426;
rommem[910] <= 16'h4A01;
rommem[911] <= 16'h6A0C;
rommem[912] <= 16'h08B9;
rommem[913] <= 16'h0001;
rommem[914] <= 16'h0001;
rommem[915] <= 16'h0427;
rommem[916] <= 16'h6000;
rommem[917] <= 16'hFEB4;
rommem[918] <= 16'h08F9;
rommem[919] <= 16'h0001;
rommem[920] <= 16'h0001;
rommem[921] <= 16'h0427;
rommem[922] <= 16'h6000;
rommem[923] <= 16'hFEA8;
rommem[924] <= 16'h2F01;
rommem[925] <= 16'h1239;
rommem[926] <= 16'h0001;
rommem[927] <= 16'h0427;
rommem[928] <= 16'h0801;
rommem[929] <= 16'h0000;
rommem[930] <= 16'h6706;
rommem[931] <= 16'h221F;
rommem[932] <= 16'h6000;
rommem[933] <= 16'hFE94;
rommem[934] <= 16'h221F;
rommem[935] <= 16'h6000;
rommem[936] <= 16'hFF12;
rommem[937] <= 16'h1239;
rommem[938] <= 16'h0001;
rommem[939] <= 16'h0426;
rommem[940] <= 16'h4239;
rommem[941] <= 16'h0001;
rommem[942] <= 16'h0426;
rommem[943] <= 16'h4A01;
rommem[944] <= 16'h6A0C;
rommem[945] <= 16'h08B9;
rommem[946] <= 16'h0000;
rommem[947] <= 16'h0001;
rommem[948] <= 16'h0427;
rommem[949] <= 16'h6000;
rommem[950] <= 16'hFE72;
rommem[951] <= 16'h08F9;
rommem[952] <= 16'h0000;
rommem[953] <= 16'h0001;
rommem[954] <= 16'h0427;
rommem[955] <= 16'h6000;
rommem[956] <= 16'hFE66;
rommem[957] <= 16'h0879;
rommem[958] <= 16'h0004;
rommem[959] <= 16'h0001;
rommem[960] <= 16'h0427;
rommem[961] <= 16'h6100;
rommem[962] <= 16'h0026;
rommem[963] <= 16'h6000;
rommem[964] <= 16'hFE56;
rommem[965] <= 16'h0879;
rommem[966] <= 16'h0005;
rommem[967] <= 16'h0001;
rommem[968] <= 16'h0427;
rommem[969] <= 16'h6100;
rommem[970] <= 16'h0016;
rommem[971] <= 16'h6000;
rommem[972] <= 16'hFE46;
rommem[973] <= 16'h0879;
rommem[974] <= 16'h0006;
rommem[975] <= 16'h0001;
rommem[976] <= 16'h0427;
rommem[977] <= 16'h6100;
rommem[978] <= 16'h0006;
rommem[979] <= 16'h6000;
rommem[980] <= 16'hFE36;
rommem[981] <= 16'h48E7;
rommem[982] <= 16'h3000;
rommem[983] <= 16'h4239;
rommem[984] <= 16'h0001;
rommem[985] <= 16'h0428;
rommem[986] <= 16'h0839;
rommem[987] <= 16'h0004;
rommem[988] <= 16'h0001;
rommem[989] <= 16'h0427;
rommem[990] <= 16'h6708;
rommem[991] <= 16'h13FC;
rommem[992] <= 16'h0002;
rommem[993] <= 16'h0001;
rommem[994] <= 16'h0428;
rommem[995] <= 16'h0839;
rommem[996] <= 16'h0005;
rommem[997] <= 16'h0001;
rommem[998] <= 16'h0427;
rommem[999] <= 16'h6708;
rommem[1000] <= 16'h08F9;
rommem[1001] <= 16'h0002;
rommem[1002] <= 16'h0001;
rommem[1003] <= 16'h0428;
rommem[1004] <= 16'h0839;
rommem[1005] <= 16'h0006;
rommem[1006] <= 16'h0001;
rommem[1007] <= 16'h0427;
rommem[1008] <= 16'h6708;
rommem[1009] <= 16'h08F9;
rommem[1010] <= 16'h0000;
rommem[1011] <= 16'h0001;
rommem[1012] <= 16'h0428;
rommem[1013] <= 16'h123C;
rommem[1014] <= 16'h00ED;
rommem[1015] <= 16'h6100;
rommem[1016] <= 16'h002C;
rommem[1017] <= 16'h6100;
rommem[1018] <= 16'hFD80;
rommem[1019] <= 16'h6100;
rommem[1020] <= 16'hFD58;
rommem[1021] <= 16'h4A01;
rommem[1022] <= 16'h6B18;
rommem[1023] <= 16'hB2BC;
rommem[1024] <= 16'h0000;
rommem[1025] <= 16'h00FA;
rommem[1026] <= 16'h1239;
rommem[1027] <= 16'h0001;
rommem[1028] <= 16'h0428;
rommem[1029] <= 16'h6100;
rommem[1030] <= 16'h0010;
rommem[1031] <= 16'h6100;
rommem[1032] <= 16'hFD64;
rommem[1033] <= 16'h6100;
rommem[1034] <= 16'hFD3C;
rommem[1035] <= 16'h4CDF;
rommem[1036] <= 16'h000C;
rommem[1037] <= 16'h4E75;
rommem[1038] <= 16'h13C1;
rommem[1039] <= 16'hFFDC;
rommem[1040] <= 16'h0000;
rommem[1041] <= 16'h4E75;
rommem[1042] <= 16'h2F03;
rommem[1043] <= 16'h263C;
rommem[1044] <= 16'h0000;
rommem[1045] <= 16'h03E8;
rommem[1046] <= 16'h51CB;
rommem[1047] <= 16'hFFFE;
rommem[1048] <= 16'h261F;
rommem[1049] <= 16'h4E75;
rommem[1050] <= 16'h2EA9;
rommem[1051] <= 16'h2EA5;
rommem[1052] <= 16'hA3A1;
rommem[1053] <= 16'hA2AC;
rommem[1054] <= 16'h2EAA;
rommem[1055] <= 16'hA8A6;
rommem[1056] <= 16'hA409;
rommem[1057] <= 16'h602E;
rommem[1058] <= 16'h2E2E;
rommem[1059] <= 16'h2E2E;
rommem[1060] <= 16'h2E71;
rommem[1061] <= 16'h312E;
rommem[1062] <= 16'h2E2E;
rommem[1063] <= 16'h7A73;
rommem[1064] <= 16'h6177;
rommem[1065] <= 16'h322E;
rommem[1066] <= 16'h2E63;
rommem[1067] <= 16'h7864;
rommem[1068] <= 16'h6534;
rommem[1069] <= 16'h332E;
rommem[1070] <= 16'h2E20;
rommem[1071] <= 16'h7666;
rommem[1072] <= 16'h7472;
rommem[1073] <= 16'h352E;
rommem[1074] <= 16'h2E6E;
rommem[1075] <= 16'h6268;
rommem[1076] <= 16'h6779;
rommem[1077] <= 16'h362E;
rommem[1078] <= 16'h2E2E;
rommem[1079] <= 16'h6D6A;
rommem[1080] <= 16'h7537;
rommem[1081] <= 16'h382E;
rommem[1082] <= 16'h2E2C;
rommem[1083] <= 16'h6B69;
rommem[1084] <= 16'h6F30;
rommem[1085] <= 16'h392E;
rommem[1086] <= 16'h2E2E;
rommem[1087] <= 16'h2F6C;
rommem[1088] <= 16'h3B70;
rommem[1089] <= 16'h2D2E;
rommem[1090] <= 16'h2E2E;
rommem[1091] <= 16'h272E;
rommem[1092] <= 16'h5B3D;
rommem[1093] <= 16'h2E2E;
rommem[1094] <= 16'hAD2E;
rommem[1095] <= 16'h0D5D;
rommem[1096] <= 16'h2E5C;
rommem[1097] <= 16'h2E2E;
rommem[1098] <= 16'h2E2E;
rommem[1099] <= 16'h2E2E;
rommem[1100] <= 16'h2E2E;
rommem[1101] <= 16'h082E;
rommem[1102] <= 16'h2E95;
rommem[1103] <= 16'h2E93;
rommem[1104] <= 16'h942E;
rommem[1105] <= 16'h2E2E;
rommem[1106] <= 16'h987F;
rommem[1107] <= 16'h922E;
rommem[1108] <= 16'h9190;
rommem[1109] <= 16'h1BAF;
rommem[1110] <= 16'hAB2E;
rommem[1111] <= 16'h972E;
rommem[1112] <= 16'h2E96;
rommem[1113] <= 16'hAE2E;
rommem[1114] <= 16'h2E2E;
rommem[1115] <= 16'h2EA7;
rommem[1116] <= 16'h2E2E;
rommem[1117] <= 16'h2E2E;
rommem[1118] <= 16'h2E2E;
rommem[1119] <= 16'h2E2E;
rommem[1120] <= 16'h2E2E;
rommem[1121] <= 16'h2E2E;
rommem[1122] <= 16'h2E2E;
rommem[1123] <= 16'h2E2E;
rommem[1124] <= 16'h2E2E;
rommem[1125] <= 16'h2E2E;
rommem[1126] <= 16'h2E2E;
rommem[1127] <= 16'h2E2E;
rommem[1128] <= 16'h2E2E;
rommem[1129] <= 16'h2E2E;
rommem[1130] <= 16'h2E2E;
rommem[1131] <= 16'h2E2E;
rommem[1132] <= 16'h2E2E;
rommem[1133] <= 16'h2E2E;
rommem[1134] <= 16'h2E2E;
rommem[1135] <= 16'h2E2E;
rommem[1136] <= 16'h2E2E;
rommem[1137] <= 16'h2E2E;
rommem[1138] <= 16'h2E2E;
rommem[1139] <= 16'h2E2E;
rommem[1140] <= 16'h2E2E;
rommem[1141] <= 16'h2E2E;
rommem[1142] <= 16'h2E2E;
rommem[1143] <= 16'h2E2E;
rommem[1144] <= 16'h2E2E;
rommem[1145] <= 16'h2E2E;
rommem[1146] <= 16'h2E2E;
rommem[1147] <= 16'h2E2E;
rommem[1148] <= 16'h2E2E;
rommem[1149] <= 16'h2E2E;
rommem[1150] <= 16'h2E2E;
rommem[1151] <= 16'h2E2E;
rommem[1152] <= 16'h2E2E;
rommem[1153] <= 16'h2E2E;
rommem[1154] <= 16'h2E2E;
rommem[1155] <= 16'h2E2E;
rommem[1156] <= 16'h2E2E;
rommem[1157] <= 16'h2E2E;
rommem[1158] <= 16'h2E2E;
rommem[1159] <= 16'h2E2E;
rommem[1160] <= 16'h2E2E;
rommem[1161] <= 16'h2E2E;
rommem[1162] <= 16'h2E2E;
rommem[1163] <= 16'h2E2E;
rommem[1164] <= 16'h2E2E;
rommem[1165] <= 16'h2E2E;
rommem[1166] <= 16'h2E2E;
rommem[1167] <= 16'h2E2E;
rommem[1168] <= 16'h2E2E;
rommem[1169] <= 16'h2E2E;
rommem[1170] <= 16'h2E2E;
rommem[1171] <= 16'h2E2E;
rommem[1172] <= 16'h2E2E;
rommem[1173] <= 16'h2E2E;
rommem[1174] <= 16'h2E2E;
rommem[1175] <= 16'hFA2E;
rommem[1176] <= 16'h2E2E;
rommem[1177] <= 16'h2E2E;
rommem[1178] <= 16'h2E2E;
rommem[1179] <= 16'h2E2E;
rommem[1180] <= 16'h2E2E;
rommem[1181] <= 16'h2E2E;
rommem[1182] <= 16'h2E2E;
rommem[1183] <= 16'h2E2E;
rommem[1184] <= 16'h2E09;
rommem[1185] <= 16'h7E2E;
rommem[1186] <= 16'h2E2E;
rommem[1187] <= 16'h2E2E;
rommem[1188] <= 16'h2E51;
rommem[1189] <= 16'h212E;
rommem[1190] <= 16'h2E2E;
rommem[1191] <= 16'h5A53;
rommem[1192] <= 16'h4157;
rommem[1193] <= 16'h402E;
rommem[1194] <= 16'h2E43;
rommem[1195] <= 16'h5844;
rommem[1196] <= 16'h4524;
rommem[1197] <= 16'h232E;
rommem[1198] <= 16'h2E20;
rommem[1199] <= 16'h5646;
rommem[1200] <= 16'h5452;
rommem[1201] <= 16'h252E;
rommem[1202] <= 16'h2E4E;
rommem[1203] <= 16'h4248;
rommem[1204] <= 16'h4759;
rommem[1205] <= 16'h5E2E;
rommem[1206] <= 16'h2E2E;
rommem[1207] <= 16'h4D4A;
rommem[1208] <= 16'h5526;
rommem[1209] <= 16'h2A2E;
rommem[1210] <= 16'h2E3C;
rommem[1211] <= 16'h4B49;
rommem[1212] <= 16'h4F29;
rommem[1213] <= 16'h282E;
rommem[1214] <= 16'h2E3E;
rommem[1215] <= 16'h3F4C;
rommem[1216] <= 16'h3A50;
rommem[1217] <= 16'h5F2E;
rommem[1218] <= 16'h2E2E;
rommem[1219] <= 16'h222E;
rommem[1220] <= 16'h7B2B;
rommem[1221] <= 16'h2E2E;
rommem[1222] <= 16'h2E2E;
rommem[1223] <= 16'h0D7D;
rommem[1224] <= 16'h2E7C;
rommem[1225] <= 16'h2E2E;
rommem[1226] <= 16'h2E2E;
rommem[1227] <= 16'h2E2E;
rommem[1228] <= 16'h2E2E;
rommem[1229] <= 16'h082E;
rommem[1230] <= 16'h2E2E;
rommem[1231] <= 16'h2E2E;
rommem[1232] <= 16'h2E2E;
rommem[1233] <= 16'h2E2E;
rommem[1234] <= 16'h2E7F;
rommem[1235] <= 16'h2E2E;
rommem[1236] <= 16'h2E2E;
rommem[1237] <= 16'h1B2E;
rommem[1238] <= 16'h2E2E;
rommem[1239] <= 16'h2E2E;
rommem[1240] <= 16'h2E2E;
rommem[1241] <= 16'h2E2E;
rommem[1242] <= 16'h2E2E;
rommem[1243] <= 16'h2E2E;
rommem[1244] <= 16'h2E2E;
rommem[1245] <= 16'h2E2E;
rommem[1246] <= 16'h2E2E;
rommem[1247] <= 16'h2E2E;
rommem[1248] <= 16'h2E2E;
rommem[1249] <= 16'h2E2E;
rommem[1250] <= 16'h2E2E;
rommem[1251] <= 16'h2E2E;
rommem[1252] <= 16'h2E2E;
rommem[1253] <= 16'h2E2E;
rommem[1254] <= 16'h2E2E;
rommem[1255] <= 16'h2E2E;
rommem[1256] <= 16'h2E2E;
rommem[1257] <= 16'h2E2E;
rommem[1258] <= 16'h2E2E;
rommem[1259] <= 16'h2E2E;
rommem[1260] <= 16'h2E2E;
rommem[1261] <= 16'h2E2E;
rommem[1262] <= 16'h2E2E;
rommem[1263] <= 16'h2E2E;
rommem[1264] <= 16'h2E2E;
rommem[1265] <= 16'h2E2E;
rommem[1266] <= 16'h2E2E;
rommem[1267] <= 16'h2E2E;
rommem[1268] <= 16'h2E2E;
rommem[1269] <= 16'h2E2E;
rommem[1270] <= 16'h2E2E;
rommem[1271] <= 16'h2E2E;
rommem[1272] <= 16'h2E2E;
rommem[1273] <= 16'h2E2E;
rommem[1274] <= 16'h2E2E;
rommem[1275] <= 16'h2E2E;
rommem[1276] <= 16'h2E2E;
rommem[1277] <= 16'h2E2E;
rommem[1278] <= 16'h2E2E;
rommem[1279] <= 16'h2E2E;
rommem[1280] <= 16'h2E2E;
rommem[1281] <= 16'h2E2E;
rommem[1282] <= 16'h2E2E;
rommem[1283] <= 16'h2E2E;
rommem[1284] <= 16'h2E2E;
rommem[1285] <= 16'h2E2E;
rommem[1286] <= 16'h2E2E;
rommem[1287] <= 16'h2E2E;
rommem[1288] <= 16'h2E2E;
rommem[1289] <= 16'h2E2E;
rommem[1290] <= 16'h2E2E;
rommem[1291] <= 16'h2E2E;
rommem[1292] <= 16'h2E2E;
rommem[1293] <= 16'h2E2E;
rommem[1294] <= 16'h2E2E;
rommem[1295] <= 16'h2E2E;
rommem[1296] <= 16'h2E2E;
rommem[1297] <= 16'h2E2E;
rommem[1298] <= 16'h2E2E;
rommem[1299] <= 16'h2E2E;
rommem[1300] <= 16'h2E2E;
rommem[1301] <= 16'h2E2E;
rommem[1302] <= 16'h2E2E;
rommem[1303] <= 16'h2E2E;
rommem[1304] <= 16'h2E2E;
rommem[1305] <= 16'h2E2E;
rommem[1306] <= 16'h2E2E;
rommem[1307] <= 16'h2E2E;
rommem[1308] <= 16'h2E2E;
rommem[1309] <= 16'h2E2E;
rommem[1310] <= 16'h2E2E;
rommem[1311] <= 16'h2E2E;
rommem[1312] <= 16'h2E09;
rommem[1313] <= 16'h7E2E;
rommem[1314] <= 16'h2E2E;
rommem[1315] <= 16'h2E2E;
rommem[1316] <= 16'h2E11;
rommem[1317] <= 16'h212E;
rommem[1318] <= 16'h2E2E;
rommem[1319] <= 16'h1A13;
rommem[1320] <= 16'h0117;
rommem[1321] <= 16'h402E;
rommem[1322] <= 16'h2E03;
rommem[1323] <= 16'h1804;
rommem[1324] <= 16'h0524;
rommem[1325] <= 16'h232E;
rommem[1326] <= 16'h2E20;
rommem[1327] <= 16'h1606;
rommem[1328] <= 16'h1412;
rommem[1329] <= 16'h252E;
rommem[1330] <= 16'h2E0E;
rommem[1331] <= 16'h0208;
rommem[1332] <= 16'h0719;
rommem[1333] <= 16'h5E2E;
rommem[1334] <= 16'h2E2E;
rommem[1335] <= 16'h0D0A;
rommem[1336] <= 16'h1526;
rommem[1337] <= 16'h2A2E;
rommem[1338] <= 16'h2E3C;
rommem[1339] <= 16'h0B09;
rommem[1340] <= 16'h0F29;
rommem[1341] <= 16'h282E;
rommem[1342] <= 16'h2E3E;
rommem[1343] <= 16'h3F0C;
rommem[1344] <= 16'h3A10;
rommem[1345] <= 16'h5F2E;
rommem[1346] <= 16'h2E2E;
rommem[1347] <= 16'h222E;
rommem[1348] <= 16'h7B2B;
rommem[1349] <= 16'h2E2E;
rommem[1350] <= 16'h2E2E;
rommem[1351] <= 16'h0D7D;
rommem[1352] <= 16'h2E7C;
rommem[1353] <= 16'h2E2E;
rommem[1354] <= 16'h2E2E;
rommem[1355] <= 16'h2E2E;
rommem[1356] <= 16'h2E2E;
rommem[1357] <= 16'h082E;
rommem[1358] <= 16'h2E2E;
rommem[1359] <= 16'h2E2E;
rommem[1360] <= 16'h2E2E;
rommem[1361] <= 16'h2E2E;
rommem[1362] <= 16'h2E7F;
rommem[1363] <= 16'h2E2E;
rommem[1364] <= 16'h2E2E;
rommem[1365] <= 16'h1B2E;
rommem[1366] <= 16'h2E2E;
rommem[1367] <= 16'h2E2E;
rommem[1368] <= 16'h2E2E;
rommem[1369] <= 16'h2E2E;
rommem[1370] <= 16'h2E2E;
rommem[1371] <= 16'h2E2E;
rommem[1372] <= 16'hA3A1;
rommem[1373] <= 16'hA22E;
rommem[1374] <= 16'h2E2E;
rommem[1375] <= 16'h2E2E;
rommem[1376] <= 16'h2E2E;
rommem[1377] <= 16'h2E2E;
rommem[1378] <= 16'h2E2E;
rommem[1379] <= 16'h2E2E;
rommem[1380] <= 16'h2E2E;
rommem[1381] <= 16'h2E2E;
rommem[1382] <= 16'h2E2E;
rommem[1383] <= 16'h2E2E;
rommem[1384] <= 16'h2E2E;
rommem[1385] <= 16'h2E2E;
rommem[1386] <= 16'h2E2E;
rommem[1387] <= 16'h2E2E;
rommem[1388] <= 16'h2E2E;
rommem[1389] <= 16'h2E2E;
rommem[1390] <= 16'h2E2E;
rommem[1391] <= 16'h2E2E;
rommem[1392] <= 16'h2E2E;
rommem[1393] <= 16'h2E2E;
rommem[1394] <= 16'h2E2E;
rommem[1395] <= 16'h2E2E;
rommem[1396] <= 16'h2E2E;
rommem[1397] <= 16'h2E2E;
rommem[1398] <= 16'h2E2E;
rommem[1399] <= 16'h2E2E;
rommem[1400] <= 16'h2E2E;
rommem[1401] <= 16'h2E2E;
rommem[1402] <= 16'h2E2E;
rommem[1403] <= 16'h2E2E;
rommem[1404] <= 16'h2E2E;
rommem[1405] <= 16'h2E2E;
rommem[1406] <= 16'h2E2E;
rommem[1407] <= 16'h2E2E;
rommem[1408] <= 16'h2E2E;
rommem[1409] <= 16'h2E2E;
rommem[1410] <= 16'h2E2E;
rommem[1411] <= 16'h2E2E;
rommem[1412] <= 16'h2E2E;
rommem[1413] <= 16'h2E2E;
rommem[1414] <= 16'h2E2E;
rommem[1415] <= 16'h2E2E;
rommem[1416] <= 16'h2E2E;
rommem[1417] <= 16'h2E2E;
rommem[1418] <= 16'h2E2E;
rommem[1419] <= 16'h2E2E;
rommem[1420] <= 16'h2E2E;
rommem[1421] <= 16'h2E2E;
rommem[1422] <= 16'h2E95;
rommem[1423] <= 16'h2E93;
rommem[1424] <= 16'h942E;
rommem[1425] <= 16'h2E2E;
rommem[1426] <= 16'h9899;
rommem[1427] <= 16'h922E;
rommem[1428] <= 16'h9190;
rommem[1429] <= 16'h2E2E;
rommem[1430] <= 16'h2E2E;
rommem[1431] <= 16'h972E;
rommem[1432] <= 16'h2E96;
rommem[1433] <= 16'h2E2E;
rommem[1434] <= 16'h4239;
rommem[1435] <= 16'h0001;
rommem[1436] <= 16'h0424;
rommem[1437] <= 16'h6100;
rommem[1438] <= 16'hF5B4;
rommem[1439] <= 16'h123C;
rommem[1440] <= 16'h0024;
rommem[1441] <= 16'h6100;
rommem[1442] <= 16'hF5F6;
rommem[1443] <= 16'h6100;
rommem[1444] <= 16'hFA66;
rommem[1445] <= 16'h0C01;
rommem[1446] <= 16'h000D;
rommem[1447] <= 16'h6706;
rommem[1448] <= 16'h6100;
rommem[1449] <= 16'hF5E8;
rommem[1450] <= 16'h60F0;
rommem[1451] <= 16'h4239;
rommem[1452] <= 16'h0001;
rommem[1453] <= 16'h0419;
rommem[1454] <= 16'h6100;
rommem[1455] <= 16'hF5AC;
rommem[1456] <= 16'h1218;
rommem[1457] <= 16'h0C01;
rommem[1458] <= 16'h0024;
rommem[1459] <= 16'h6602;
rommem[1460] <= 16'h1218;
rommem[1461] <= 16'h0C01;
rommem[1462] <= 16'h0067;
rommem[1463] <= 16'h6700;
rommem[1464] <= 16'h0640;
rommem[1465] <= 16'h0C01;
rommem[1466] <= 16'h003A;
rommem[1467] <= 16'h6700;
rommem[1468] <= 16'h0156;
rommem[1469] <= 16'h0C01;
rommem[1470] <= 16'h0044;
rommem[1471] <= 16'h6700;
rommem[1472] <= 16'h01BC;
rommem[1473] <= 16'h0C01;
rommem[1474] <= 16'h0046;
rommem[1475] <= 16'h6700;
rommem[1476] <= 16'h00F0;
rommem[1477] <= 16'h0C01;
rommem[1478] <= 16'h0042;
rommem[1479] <= 16'h6700;
rommem[1480] <= 16'hFFFF;
rommem[1481] <= 16'h0C01;
rommem[1482] <= 16'h004A;
rommem[1483] <= 16'h6700;
rommem[1484] <= 16'h0194;
rommem[1485] <= 16'h0C01;
rommem[1486] <= 16'h004C;
rommem[1487] <= 16'h6700;
rommem[1488] <= 16'h0328;
rommem[1489] <= 16'h0C01;
rommem[1490] <= 16'h003F;
rommem[1491] <= 16'h6724;
rommem[1492] <= 16'h0C01;
rommem[1493] <= 16'h0043;
rommem[1494] <= 16'h6702;
rommem[1495] <= 16'h6084;
rommem[1496] <= 16'h1218;
rommem[1497] <= 16'h0C01;
rommem[1498] <= 16'h004C;
rommem[1499] <= 16'h6600;
rommem[1500] <= 16'hFF7C;
rommem[1501] <= 16'h1218;
rommem[1502] <= 16'h0C01;
rommem[1503] <= 16'h0053;
rommem[1504] <= 16'h6600;
rommem[1505] <= 16'hFF72;
rommem[1506] <= 16'h6100;
rommem[1507] <= 16'h0216;
rommem[1508] <= 16'h6000;
rommem[1509] <= 16'hFF6A;
rommem[1510] <= 16'h43F9;
rommem[1511] <= 16'hFFFC;
rommem[1512] <= 16'h0BDC;
rommem[1513] <= 16'h4EB9;
rommem[1514] <= 16'hFFFC;
rommem[1515] <= 16'h02AA;
rommem[1516] <= 16'h6000;
rommem[1517] <= 16'hFF5A;
rommem[1518] <= 16'h3F20;
rommem[1519] <= 16'h3D20;
rommem[1520] <= 16'h4469;
rommem[1521] <= 16'h7370;
rommem[1522] <= 16'h6C61;
rommem[1523] <= 16'h7920;
rommem[1524] <= 16'h6865;
rommem[1525] <= 16'h6C70;
rommem[1526] <= 16'h0D0A;
rommem[1527] <= 16'h434C;
rommem[1528] <= 16'h5320;
rommem[1529] <= 16'h3D20;
rommem[1530] <= 16'h636C;
rommem[1531] <= 16'h6561;
rommem[1532] <= 16'h7220;
rommem[1533] <= 16'h7363;
rommem[1534] <= 16'h7265;
rommem[1535] <= 16'h656E;
rommem[1536] <= 16'h0D0A;
rommem[1537] <= 16'h3A20;
rommem[1538] <= 16'h3D20;
rommem[1539] <= 16'h4564;
rommem[1540] <= 16'h6974;
rommem[1541] <= 16'h206D;
rommem[1542] <= 16'h656D;
rommem[1543] <= 16'h6F72;
rommem[1544] <= 16'h7920;
rommem[1545] <= 16'h6279;
rommem[1546] <= 16'h7465;
rommem[1547] <= 16'h730D;
rommem[1548] <= 16'h0A46;
rommem[1549] <= 16'h203D;
rommem[1550] <= 16'h2046;
rommem[1551] <= 16'h696C;
rommem[1552] <= 16'h6C20;
rommem[1553] <= 16'h6D65;
rommem[1554] <= 16'h6D6F;
rommem[1555] <= 16'h7279;
rommem[1556] <= 16'h0D0A;
rommem[1557] <= 16'h4C20;
rommem[1558] <= 16'h3D20;
rommem[1559] <= 16'h4C6F;
rommem[1560] <= 16'h6164;
rommem[1561] <= 16'h2053;
rommem[1562] <= 16'h3139;
rommem[1563] <= 16'h2066;
rommem[1564] <= 16'h696C;
rommem[1565] <= 16'h650D;
rommem[1566] <= 16'h0A44;
rommem[1567] <= 16'h203D;
rommem[1568] <= 16'h2044;
rommem[1569] <= 16'h756D;
rommem[1570] <= 16'h7020;
rommem[1571] <= 16'h6D65;
rommem[1572] <= 16'h6D6F;
rommem[1573] <= 16'h7279;
rommem[1574] <= 16'h0D0A;
rommem[1575] <= 16'h4220;
rommem[1576] <= 16'h3D20;
rommem[1577] <= 16'h7374;
rommem[1578] <= 16'h6172;
rommem[1579] <= 16'h7420;
rommem[1580] <= 16'h7469;
rommem[1581] <= 16'h6E79;
rommem[1582] <= 16'h2062;
rommem[1583] <= 16'h6173;
rommem[1584] <= 16'h6963;
rommem[1585] <= 16'h0D0A;
rommem[1586] <= 16'h4A20;
rommem[1587] <= 16'h3D20;
rommem[1588] <= 16'h4A75;
rommem[1589] <= 16'h6D70;
rommem[1590] <= 16'h2074;
rommem[1591] <= 16'h6F20;
rommem[1592] <= 16'h636F;
rommem[1593] <= 16'h6465;
rommem[1594] <= 16'h0D0A;
rommem[1595] <= 16'h00FF;
rommem[1596] <= 16'h1218;
rommem[1597] <= 16'h1801;
rommem[1598] <= 16'h6100;
rommem[1599] <= 16'h0044;
rommem[1600] <= 16'h6100;
rommem[1601] <= 16'h00EE;
rommem[1602] <= 16'h2241;
rommem[1603] <= 16'h6100;
rommem[1604] <= 16'h003A;
rommem[1605] <= 16'h6100;
rommem[1606] <= 16'h00E4;
rommem[1607] <= 16'h2601;
rommem[1608] <= 16'h6100;
rommem[1609] <= 16'h0030;
rommem[1610] <= 16'h6100;
rommem[1611] <= 16'h00DA;
rommem[1612] <= 16'h0C04;
rommem[1613] <= 16'h004C;
rommem[1614] <= 16'h660A;
rommem[1615] <= 16'h22C1;
rommem[1616] <= 16'h51CB;
rommem[1617] <= 16'hFFFC;
rommem[1618] <= 16'h6000;
rommem[1619] <= 16'hFE8E;
rommem[1620] <= 16'h0C04;
rommem[1621] <= 16'h0057;
rommem[1622] <= 16'h660A;
rommem[1623] <= 16'h32C1;
rommem[1624] <= 16'h51CB;
rommem[1625] <= 16'hFFFC;
rommem[1626] <= 16'h6000;
rommem[1627] <= 16'hFE7E;
rommem[1628] <= 16'h12C1;
rommem[1629] <= 16'h51CB;
rommem[1630] <= 16'hFFFC;
rommem[1631] <= 16'h6000;
rommem[1632] <= 16'hFE74;
rommem[1633] <= 16'h1218;
rommem[1634] <= 16'h0C01;
rommem[1635] <= 16'h0020;
rommem[1636] <= 16'h67F8;
rommem[1637] <= 16'h5388;
rommem[1638] <= 16'h4E75;
rommem[1639] <= 16'h6100;
rommem[1640] <= 16'hFFF2;
rommem[1641] <= 16'h6100;
rommem[1642] <= 16'h009C;
rommem[1643] <= 16'h2241;
rommem[1644] <= 16'h6100;
rommem[1645] <= 16'hFFE8;
rommem[1646] <= 16'h6100;
rommem[1647] <= 16'h0092;
rommem[1648] <= 16'h12C1;
rommem[1649] <= 16'h6100;
rommem[1650] <= 16'hFFDE;
rommem[1651] <= 16'h6100;
rommem[1652] <= 16'h0088;
rommem[1653] <= 16'h12C1;
rommem[1654] <= 16'h6100;
rommem[1655] <= 16'hFFD4;
rommem[1656] <= 16'h6100;
rommem[1657] <= 16'h007E;
rommem[1658] <= 16'h12C1;
rommem[1659] <= 16'h6100;
rommem[1660] <= 16'hFFCA;
rommem[1661] <= 16'h6100;
rommem[1662] <= 16'h0074;
rommem[1663] <= 16'h12C1;
rommem[1664] <= 16'h6100;
rommem[1665] <= 16'hFFC0;
rommem[1666] <= 16'h6100;
rommem[1667] <= 16'h006A;
rommem[1668] <= 16'h12C1;
rommem[1669] <= 16'h6100;
rommem[1670] <= 16'hFFB6;
rommem[1671] <= 16'h6100;
rommem[1672] <= 16'h0060;
rommem[1673] <= 16'h12C1;
rommem[1674] <= 16'h6100;
rommem[1675] <= 16'hFFAC;
rommem[1676] <= 16'h6100;
rommem[1677] <= 16'h0056;
rommem[1678] <= 16'h12C1;
rommem[1679] <= 16'h6100;
rommem[1680] <= 16'hFFA2;
rommem[1681] <= 16'h6100;
rommem[1682] <= 16'h004C;
rommem[1683] <= 16'h12C1;
rommem[1684] <= 16'h6000;
rommem[1685] <= 16'hFE0A;
rommem[1686] <= 16'h6100;
rommem[1687] <= 16'hFF94;
rommem[1688] <= 16'h6100;
rommem[1689] <= 16'h003E;
rommem[1690] <= 16'h2041;
rommem[1691] <= 16'h4E90;
rommem[1692] <= 16'h6000;
rommem[1693] <= 16'hFDFA;
rommem[1694] <= 16'h6100;
rommem[1695] <= 16'hFF84;
rommem[1696] <= 16'h6100;
rommem[1697] <= 16'h002E;
rommem[1698] <= 16'h2041;
rommem[1699] <= 16'h4EB9;
rommem[1700] <= 16'hFFFC;
rommem[1701] <= 16'h00F0;
rommem[1702] <= 16'h6100;
rommem[1703] <= 16'hF7B8;
rommem[1704] <= 16'h6100;
rommem[1705] <= 16'hF7B4;
rommem[1706] <= 16'h6100;
rommem[1707] <= 16'hF7B0;
rommem[1708] <= 16'h6100;
rommem[1709] <= 16'hF7AC;
rommem[1710] <= 16'h6100;
rommem[1711] <= 16'hF7A8;
rommem[1712] <= 16'h6100;
rommem[1713] <= 16'hF7A4;
rommem[1714] <= 16'h6100;
rommem[1715] <= 16'hF7A0;
rommem[1716] <= 16'h6100;
rommem[1717] <= 16'hF79C;
rommem[1718] <= 16'h6000;
rommem[1719] <= 16'hFDC6;
rommem[1720] <= 16'h48E7;
rommem[1721] <= 16'hA000;
rommem[1722] <= 16'h4282;
rommem[1723] <= 16'h7007;
rommem[1724] <= 16'h1218;
rommem[1725] <= 16'h6100;
rommem[1726] <= 16'h001E;
rommem[1727] <= 16'hB23C;
rommem[1728] <= 16'h00FF;
rommem[1729] <= 16'h670E;
rommem[1730] <= 16'hE98A;
rommem[1731] <= 16'h0281;
rommem[1732] <= 16'h0000;
rommem[1733] <= 16'h000F;
rommem[1734] <= 16'h8481;
rommem[1735] <= 16'h51C8;
rommem[1736] <= 16'hFFE8;
rommem[1737] <= 16'h2202;
rommem[1738] <= 16'h4CDF;
rommem[1739] <= 16'h0005;
rommem[1740] <= 16'h4E75;
rommem[1741] <= 16'h0C01;
rommem[1742] <= 16'h0030;
rommem[1743] <= 16'h6538;
rommem[1744] <= 16'h0C01;
rommem[1745] <= 16'h0039;
rommem[1746] <= 16'h6206;
rommem[1747] <= 16'h0401;
rommem[1748] <= 16'h0030;
rommem[1749] <= 16'h4E75;
rommem[1750] <= 16'h0C01;
rommem[1751] <= 16'h0041;
rommem[1752] <= 16'h6526;
rommem[1753] <= 16'h0C01;
rommem[1754] <= 16'h0046;
rommem[1755] <= 16'h620A;
rommem[1756] <= 16'h0401;
rommem[1757] <= 16'h0041;
rommem[1758] <= 16'h0601;
rommem[1759] <= 16'h000A;
rommem[1760] <= 16'h4E75;
rommem[1761] <= 16'h0C01;
rommem[1762] <= 16'h0061;
rommem[1763] <= 16'h6510;
rommem[1764] <= 16'h0C01;
rommem[1765] <= 16'h0066;
rommem[1766] <= 16'h620A;
rommem[1767] <= 16'h0401;
rommem[1768] <= 16'h0061;
rommem[1769] <= 16'h0601;
rommem[1770] <= 16'h000A;
rommem[1771] <= 16'h4E75;
rommem[1772] <= 16'h72FF;
rommem[1773] <= 16'h4E75;
rommem[1774] <= 16'h4BF9;
rommem[1775] <= 16'hFFE0;
rommem[1776] <= 16'h0000;
rommem[1777] <= 16'h302D;
rommem[1778] <= 16'h04AC;
rommem[1779] <= 16'h0800;
rommem[1780] <= 16'h000D;
rommem[1781] <= 16'h67F6;
rommem[1782] <= 16'h2B7C;
rommem[1783] <= 16'h0001;
rommem[1784] <= 16'h4000;
rommem[1785] <= 16'h04BC;
rommem[1786] <= 16'h3B79;
rommem[1787] <= 16'h0001;
rommem[1788] <= 16'h0004;
rommem[1789] <= 16'h04A8;
rommem[1790] <= 16'h2B7C;
rommem[1791] <= 16'h0000;
rommem[1792] <= 16'h0000;
rommem[1793] <= 16'h0498;
rommem[1794] <= 16'h2B7C;
rommem[1795] <= 16'h0000;
rommem[1796] <= 16'h0140;
rommem[1797] <= 16'h04A4;
rommem[1798] <= 16'h2B7C;
rommem[1799] <= 16'h0000;
rommem[1800] <= 16'h0000;
rommem[1801] <= 16'h049C;
rommem[1802] <= 16'h3B7C;
rommem[1803] <= 16'h8080;
rommem[1804] <= 16'h04AC;
rommem[1805] <= 16'h4E75;
rommem[1806] <= 16'h48E7;
rommem[1807] <= 16'h8004;
rommem[1808] <= 16'h4BF9;
rommem[1809] <= 16'hFFE0;
rommem[1810] <= 16'h0000;
rommem[1811] <= 16'h302D;
rommem[1812] <= 16'h04AC;
rommem[1813] <= 16'h0800;
rommem[1814] <= 16'h000D;
rommem[1815] <= 16'h67F6;
rommem[1816] <= 16'h2B7C;
rommem[1817] <= 16'h0001;
rommem[1818] <= 16'h3600;
rommem[1819] <= 16'h04B0;
rommem[1820] <= 16'h2B7C;
rommem[1821] <= 16'h0000;
rommem[1822] <= 16'h0A00;
rommem[1823] <= 16'h0480;
rommem[1824] <= 16'h2B7C;
rommem[1825] <= 16'h0000;
rommem[1826] <= 16'h0000;
rommem[1827] <= 16'h0484;
rommem[1828] <= 16'h2B7C;
rommem[1829] <= 16'h0001;
rommem[1830] <= 16'h3600;
rommem[1831] <= 16'h04BC;
rommem[1832] <= 16'h2B7C;
rommem[1833] <= 16'h0000;
rommem[1834] <= 16'h0000;
rommem[1835] <= 16'h0498;
rommem[1836] <= 16'h2B7C;
rommem[1837] <= 16'h0000;
rommem[1838] <= 16'h0000;
rommem[1839] <= 16'h049C;
rommem[1840] <= 16'h2B7C;
rommem[1841] <= 16'hFFFF;
rommem[1842] <= 16'hFFFF;
rommem[1843] <= 16'h04A0;
rommem[1844] <= 16'h2B7C;
rommem[1845] <= 16'hFFFF;
rommem[1846] <= 16'hFFFF;
rommem[1847] <= 16'h04A4;
rommem[1848] <= 16'h3B7C;
rommem[1849] <= 16'h0011;
rommem[1850] <= 16'h04AE;
rommem[1851] <= 16'h3B7C;
rommem[1852] <= 16'h8082;
rommem[1853] <= 16'h04AC;
rommem[1854] <= 16'h4CDF;
rommem[1855] <= 16'h2001;
rommem[1856] <= 16'h48E7;
rommem[1857] <= 16'h8004;
rommem[1858] <= 16'h4BF9;
rommem[1859] <= 16'hFFE0;
rommem[1860] <= 16'h0000;
rommem[1861] <= 16'h302D;
rommem[1862] <= 16'h04AC;
rommem[1863] <= 16'h0800;
rommem[1864] <= 16'h000D;
rommem[1865] <= 16'h67F6;
rommem[1866] <= 16'h2B7C;
rommem[1867] <= 16'h0000;
rommem[1868] <= 16'h0A00;
rommem[1869] <= 16'h04BC;
rommem[1870] <= 16'h2B7C;
rommem[1871] <= 16'h0001;
rommem[1872] <= 16'h3600;
rommem[1873] <= 16'h0498;
rommem[1874] <= 16'h2B7C;
rommem[1875] <= 16'h0000;
rommem[1876] <= 16'h0000;
rommem[1877] <= 16'h049C;
rommem[1878] <= 16'h2B7C;
rommem[1879] <= 16'hFFFF;
rommem[1880] <= 16'hFFFF;
rommem[1881] <= 16'h04A4;
rommem[1882] <= 16'h3B79;
rommem[1883] <= 16'h0001;
rommem[1884] <= 16'h0004;
rommem[1885] <= 16'h04A8;
rommem[1886] <= 16'h3B7C;
rommem[1887] <= 16'h8080;
rommem[1888] <= 16'h04AC;
rommem[1889] <= 16'h4CDF;
rommem[1890] <= 16'h2001;
rommem[1891] <= 16'h4E75;
rommem[1892] <= 16'h600A;
rommem[1893] <= 16'h6100;
rommem[1894] <= 16'h017A;
rommem[1895] <= 16'h0C00;
rommem[1896] <= 16'h000A;
rommem[1897] <= 16'h66F6;
rommem[1898] <= 16'h6100;
rommem[1899] <= 16'h0170;
rommem[1900] <= 16'h1800;
rommem[1901] <= 16'h0C04;
rommem[1902] <= 16'h001A;
rommem[1903] <= 16'h6700;
rommem[1904] <= 16'hFC54;
rommem[1905] <= 16'h0C04;
rommem[1906] <= 16'h0053;
rommem[1907] <= 16'h66E2;
rommem[1908] <= 16'h6100;
rommem[1909] <= 16'h015C;
rommem[1910] <= 16'h1800;
rommem[1911] <= 16'h0C04;
rommem[1912] <= 16'h0030;
rommem[1913] <= 16'h65D6;
rommem[1914] <= 16'h0C04;
rommem[1915] <= 16'h0039;
rommem[1916] <= 16'h62D0;
rommem[1917] <= 16'h6100;
rommem[1918] <= 16'h014A;
rommem[1919] <= 16'h6100;
rommem[1920] <= 16'hFE9A;
rommem[1921] <= 16'h1401;
rommem[1922] <= 16'h6100;
rommem[1923] <= 16'h0140;
rommem[1924] <= 16'h6100;
rommem[1925] <= 16'hFE90;
rommem[1926] <= 16'hE90A;
rommem[1927] <= 16'h8202;
rommem[1928] <= 16'h1601;
rommem[1929] <= 16'h0C04;
rommem[1930] <= 16'h0030;
rommem[1931] <= 16'h67B2;
rommem[1932] <= 16'h0C04;
rommem[1933] <= 16'h0031;
rommem[1934] <= 16'h676A;
rommem[1935] <= 16'h0C04;
rommem[1936] <= 16'h0032;
rommem[1937] <= 16'h676A;
rommem[1938] <= 16'h0C04;
rommem[1939] <= 16'h0033;
rommem[1940] <= 16'h676A;
rommem[1941] <= 16'h0C04;
rommem[1942] <= 16'h0035;
rommem[1943] <= 16'h679A;
rommem[1944] <= 16'h0C04;
rommem[1945] <= 16'h0037;
rommem[1946] <= 16'h6764;
rommem[1947] <= 16'h0C04;
rommem[1948] <= 16'h0038;
rommem[1949] <= 16'h676C;
rommem[1950] <= 16'h0C04;
rommem[1951] <= 16'h0039;
rommem[1952] <= 16'h6774;
rommem[1953] <= 16'h6086;
rommem[1954] <= 16'h0243;
rommem[1955] <= 16'h00FF;
rommem[1956] <= 16'h5343;
rommem[1957] <= 16'h4282;
rommem[1958] <= 16'h6100;
rommem[1959] <= 16'h00F8;
rommem[1960] <= 16'h6100;
rommem[1961] <= 16'hFE48;
rommem[1962] <= 16'hE98A;
rommem[1963] <= 16'h8401;
rommem[1964] <= 16'h6100;
rommem[1965] <= 16'h00EC;
rommem[1966] <= 16'h6100;
rommem[1967] <= 16'hFE3C;
rommem[1968] <= 16'hE98A;
rommem[1969] <= 16'h8401;
rommem[1970] <= 16'h12C2;
rommem[1971] <= 16'h51CB;
rommem[1972] <= 16'hFFE2;
rommem[1973] <= 16'h4282;
rommem[1974] <= 16'h6100;
rommem[1975] <= 16'h00D8;
rommem[1976] <= 16'h6100;
rommem[1977] <= 16'hFE28;
rommem[1978] <= 16'hE98A;
rommem[1979] <= 16'h8401;
rommem[1980] <= 16'h6100;
rommem[1981] <= 16'h00CC;
rommem[1982] <= 16'h6100;
rommem[1983] <= 16'hFE1C;
rommem[1984] <= 16'hE98A;
rommem[1985] <= 16'h8401;
rommem[1986] <= 16'h6000;
rommem[1987] <= 16'hFF44;
rommem[1988] <= 16'h6100;
rommem[1989] <= 16'h003A;
rommem[1990] <= 16'h60B6;
rommem[1991] <= 16'h6100;
rommem[1992] <= 16'h0042;
rommem[1993] <= 16'h60B0;
rommem[1994] <= 16'h6100;
rommem[1995] <= 16'h004A;
rommem[1996] <= 16'h60AA;
rommem[1997] <= 16'h6100;
rommem[1998] <= 16'h0044;
rommem[1999] <= 16'h23C9;
rommem[2000] <= 16'h0000;
rommem[2001] <= 16'h0000;
rommem[2002] <= 16'h6000;
rommem[2003] <= 16'hFB8E;
rommem[2004] <= 16'h6100;
rommem[2005] <= 16'h0028;
rommem[2006] <= 16'h23C9;
rommem[2007] <= 16'h0000;
rommem[2008] <= 16'h0000;
rommem[2009] <= 16'h6000;
rommem[2010] <= 16'hFB80;
rommem[2011] <= 16'h6100;
rommem[2012] <= 16'h000C;
rommem[2013] <= 16'h23C9;
rommem[2014] <= 16'h0000;
rommem[2015] <= 16'h0000;
rommem[2016] <= 16'h6000;
rommem[2017] <= 16'hFB72;
rommem[2018] <= 16'h4282;
rommem[2019] <= 16'h6100;
rommem[2020] <= 16'h007E;
rommem[2021] <= 16'h6100;
rommem[2022] <= 16'hFDCE;
rommem[2023] <= 16'h1401;
rommem[2024] <= 16'h604A;
rommem[2025] <= 16'h4282;
rommem[2026] <= 16'h6100;
rommem[2027] <= 16'h0070;
rommem[2028] <= 16'h6100;
rommem[2029] <= 16'hFDC0;
rommem[2030] <= 16'h1401;
rommem[2031] <= 16'h6024;
rommem[2032] <= 16'h4282;
rommem[2033] <= 16'h6100;
rommem[2034] <= 16'h0062;
rommem[2035] <= 16'h6100;
rommem[2036] <= 16'hFDB2;
rommem[2037] <= 16'h1401;
rommem[2038] <= 16'h6100;
rommem[2039] <= 16'h0058;
rommem[2040] <= 16'h6100;
rommem[2041] <= 16'hFDA8;
rommem[2042] <= 16'hE98A;
rommem[2043] <= 16'h8401;
rommem[2044] <= 16'h6100;
rommem[2045] <= 16'h004C;
rommem[2046] <= 16'h6100;
rommem[2047] <= 16'hFD9C;
rommem[2048] <= 16'hE98A;
rommem[2049] <= 16'h8401;
rommem[2050] <= 16'h6100;
rommem[2051] <= 16'h0040;
rommem[2052] <= 16'h6100;
rommem[2053] <= 16'hFD90;
rommem[2054] <= 16'hE98A;
rommem[2055] <= 16'h8401;
rommem[2056] <= 16'h6100;
rommem[2057] <= 16'h0034;
rommem[2058] <= 16'h6100;
rommem[2059] <= 16'hFD84;
rommem[2060] <= 16'hE98A;
rommem[2061] <= 16'h8401;
rommem[2062] <= 16'h6100;
rommem[2063] <= 16'h0028;
rommem[2064] <= 16'h6100;
rommem[2065] <= 16'hFD78;
rommem[2066] <= 16'hE98A;
rommem[2067] <= 16'h8401;
rommem[2068] <= 16'h6100;
rommem[2069] <= 16'h001C;
rommem[2070] <= 16'h6100;
rommem[2071] <= 16'hFD6C;
rommem[2072] <= 16'hE98A;
rommem[2073] <= 16'h8401;
rommem[2074] <= 16'h6100;
rommem[2075] <= 16'h0010;
rommem[2076] <= 16'h6100;
rommem[2077] <= 16'hFD60;
rommem[2078] <= 16'hE98A;
rommem[2079] <= 16'h8401;
rommem[2080] <= 16'h4284;
rommem[2081] <= 16'h2242;
rommem[2082] <= 16'h4E75;
rommem[2083] <= 16'h6100;
rommem[2084] <= 16'hF554;
rommem[2085] <= 16'h670C;
rommem[2086] <= 16'h6100;
rommem[2087] <= 16'hF560;
rommem[2088] <= 16'h0C01;
rommem[2089] <= 16'h0000;
rommem[2090] <= 16'h6700;
rommem[2091] <= 16'hFADE;
rommem[2092] <= 16'h6100;
rommem[2093] <= 16'hFFFF;
rommem[2094] <= 16'h67E8;
rommem[2095] <= 16'h1200;
rommem[2096] <= 16'h4E75;
rommem[2097] <= 16'h33FC;
rommem[2098] <= 16'hA6A6;
rommem[2099] <= 16'hFFDC;
rommem[2100] <= 16'h0600;
rommem[2101] <= 16'h2C7C;
rommem[2102] <= 16'hFFE0;
rommem[2103] <= 16'h0000;
rommem[2104] <= 16'h343C;
rommem[2105] <= 16'h0007;
rommem[2106] <= 16'h1001;
rommem[2107] <= 16'h0240;
rommem[2108] <= 16'h000F;
rommem[2109] <= 16'h0C40;
rommem[2110] <= 16'h0009;
rommem[2111] <= 16'h6302;
rommem[2112] <= 16'h5E40;
rommem[2113] <= 16'h0640;
rommem[2114] <= 16'h0030;
rommem[2115] <= 16'h3602;
rommem[2116] <= 16'hE743;
rommem[2117] <= 16'h382E;
rommem[2118] <= 16'h042C;
rommem[2119] <= 16'hB87C;
rommem[2120] <= 16'h001C;
rommem[2121] <= 16'h64F6;
rommem[2122] <= 16'h4880;
rommem[2123] <= 16'h3D40;
rommem[2124] <= 16'h0420;
rommem[2125] <= 16'h3D7C;
rommem[2126] <= 16'h7FFF;
rommem[2127] <= 16'h0422;
rommem[2128] <= 16'h3D7C;
rommem[2129] <= 16'h000F;
rommem[2130] <= 16'h0424;
rommem[2131] <= 16'h3D43;
rommem[2132] <= 16'h0426;
rommem[2133] <= 16'h3D7C;
rommem[2134] <= 16'h0008;
rommem[2135] <= 16'h0428;
rommem[2136] <= 16'h3D7C;
rommem[2137] <= 16'h0707;
rommem[2138] <= 16'h042A;
rommem[2139] <= 16'h3D7C;
rommem[2140] <= 16'h0000;
rommem[2141] <= 16'h042E;
rommem[2142] <= 16'hE899;
rommem[2143] <= 16'h57CA;
rommem[2144] <= 16'hFFB4;
rommem[2145] <= 16'h4ED5;
rommem[2146] <= 16'h33FC;
rommem[2147] <= 16'hA5A5;
rommem[2148] <= 16'hFFDC;
rommem[2149] <= 16'h0600;
rommem[2150] <= 16'h207C;
rommem[2151] <= 16'h0003;
rommem[2152] <= 16'h0000;
rommem[2153] <= 16'h203C;
rommem[2154] <= 16'hAAAA;
rommem[2155] <= 16'h5555;
rommem[2156] <= 16'h20C0;
rommem[2157] <= 16'h2208;
rommem[2158] <= 16'h4A41;
rommem[2159] <= 16'h660A;
rommem[2160] <= 16'h4BF9;
rommem[2161] <= 16'hFFFC;
rommem[2162] <= 16'h10EA;
rommem[2163] <= 16'h6000;
rommem[2164] <= 16'hFF7A;
rommem[2165] <= 16'h33FC;
rommem[2166] <= 16'hA9A9;
rommem[2167] <= 16'hFFDC;
rommem[2168] <= 16'h0600;
rommem[2169] <= 16'hB1FC;
rommem[2170] <= 16'h0005;
rommem[2171] <= 16'hFFFC;
rommem[2172] <= 16'h66DE;
rommem[2173] <= 16'h7200;
rommem[2174] <= 16'h6100;
rommem[2175] <= 16'hF00C;
rommem[2176] <= 16'h6000;
rommem[2177] <= 16'hFC42;
rommem[2178] <= 16'h33FC;
rommem[2179] <= 16'hA7A7;
rommem[2180] <= 16'hFFDC;
rommem[2181] <= 16'h0600;
rommem[2182] <= 16'h2448;
rommem[2183] <= 16'h207C;
rommem[2184] <= 16'h0003;
rommem[2185] <= 16'h0000;
rommem[2186] <= 16'h2A18;
rommem[2187] <= 16'hB5C8;
rommem[2188] <= 16'h671A;
rommem[2189] <= 16'h2208;
rommem[2190] <= 16'h4A41;
rommem[2191] <= 16'h660A;
rommem[2192] <= 16'h4BF9;
rommem[2193] <= 16'hFFFC;
rommem[2194] <= 16'h112A;
rommem[2195] <= 16'h6000;
rommem[2196] <= 16'hFF3A;
rommem[2197] <= 16'h0C85;
rommem[2198] <= 16'hAAAA;
rommem[2199] <= 16'h5555;
rommem[2200] <= 16'h67E2;
rommem[2201] <= 16'h6678;
rommem[2202] <= 16'h33FC;
rommem[2203] <= 16'hA8A8;
rommem[2204] <= 16'hFFDC;
rommem[2205] <= 16'h0600;
rommem[2206] <= 16'h207C;
rommem[2207] <= 16'h0003;
rommem[2208] <= 16'h0000;
rommem[2209] <= 16'h203C;
rommem[2210] <= 16'h5555;
rommem[2211] <= 16'hAAAA;
rommem[2212] <= 16'h20C0;
rommem[2213] <= 16'h2208;
rommem[2214] <= 16'h4A41;
rommem[2215] <= 16'h660A;
rommem[2216] <= 16'h4BF9;
rommem[2217] <= 16'hFFFC;
rommem[2218] <= 16'h115A;
rommem[2219] <= 16'h6000;
rommem[2220] <= 16'hFF0A;
rommem[2221] <= 16'hB1FC;
rommem[2222] <= 16'h1FFF;
rommem[2223] <= 16'hFFFC;
rommem[2224] <= 16'h66E6;
rommem[2225] <= 16'h2448;
rommem[2226] <= 16'h207C;
rommem[2227] <= 16'h0003;
rommem[2228] <= 16'h0000;
rommem[2229] <= 16'h2018;
rommem[2230] <= 16'hB5C8;
rommem[2231] <= 16'h671A;
rommem[2232] <= 16'h2208;
rommem[2233] <= 16'h4A41;
rommem[2234] <= 16'h660A;
rommem[2235] <= 16'h4BF9;
rommem[2236] <= 16'hFFFC;
rommem[2237] <= 16'h1180;
rommem[2238] <= 16'h6000;
rommem[2239] <= 16'hFEE4;
rommem[2240] <= 16'h0C80;
rommem[2241] <= 16'h5555;
rommem[2242] <= 16'hAAAA;
rommem[2243] <= 16'h67E2;
rommem[2244] <= 16'h6622;
rommem[2245] <= 16'h23C8;
rommem[2246] <= 16'h0001;
rommem[2247] <= 16'h0008;
rommem[2248] <= 16'h91FC;
rommem[2249] <= 16'h0000;
rommem[2250] <= 16'h000C;
rommem[2251] <= 16'h21C8;
rommem[2252] <= 16'h0404;
rommem[2253] <= 16'h21FC;
rommem[2254] <= 16'h4652;
rommem[2255] <= 16'h4545;
rommem[2256] <= 16'h0400;
rommem[2257] <= 16'h21FC;
rommem[2258] <= 16'h0000;
rommem[2259] <= 16'h0408;
rommem[2260] <= 16'h0408;
rommem[2261] <= 16'h4ED3;
rommem[2262] <= 16'h4ED3;
rommem[2263] <= 16'h60FC;
rommem[2264] <= 16'h6100;
rommem[2265] <= 16'h0080;
rommem[2266] <= 16'h6100;
rommem[2267] <= 16'h0006;
rommem[2268] <= 16'h6000;
rommem[2269] <= 16'hF97A;
rommem[2270] <= 16'h4DF9;
rommem[2271] <= 16'hFFDC;
rommem[2272] <= 16'h0000;
rommem[2273] <= 16'h4BF9;
rommem[2274] <= 16'hFFE0;
rommem[2275] <= 16'h0000;
rommem[2276] <= 16'h2C3C;
rommem[2277] <= 16'h0003;
rommem[2278] <= 16'h0D40;
rommem[2279] <= 16'h202E;
rommem[2280] <= 16'h0C00;
rommem[2281] <= 16'h3200;
rommem[2282] <= 16'h4840;
rommem[2283] <= 16'h0240;
rommem[2284] <= 16'h00FF;
rommem[2285] <= 16'h0241;
rommem[2286] <= 16'h00FF;
rommem[2287] <= 16'h426E;
rommem[2288] <= 16'h0C04;
rommem[2289] <= 16'h242E;
rommem[2290] <= 16'h0C00;
rommem[2291] <= 16'h3602;
rommem[2292] <= 16'h4842;
rommem[2293] <= 16'h0242;
rommem[2294] <= 16'h00FF;
rommem[2295] <= 16'h0243;
rommem[2296] <= 16'h00FF;
rommem[2297] <= 16'h426E;
rommem[2298] <= 16'h0C04;
rommem[2299] <= 16'h282E;
rommem[2300] <= 16'h0C00;
rommem[2301] <= 16'h0244;
rommem[2302] <= 16'h7FFF;
rommem[2303] <= 16'h426E;
rommem[2304] <= 16'h0C04;
rommem[2305] <= 16'h3E2D;
rommem[2306] <= 16'h042C;
rommem[2307] <= 16'hBE7C;
rommem[2308] <= 16'h001C;
rommem[2309] <= 16'h64F6;
rommem[2310] <= 16'h3B7C;
rommem[2311] <= 16'h0001;
rommem[2312] <= 16'h0422;
rommem[2313] <= 16'h3B44;
rommem[2314] <= 16'h0424;
rommem[2315] <= 16'h3B40;
rommem[2316] <= 16'h0426;
rommem[2317] <= 16'h3B41;
rommem[2318] <= 16'h0428;
rommem[2319] <= 16'h3B42;
rommem[2320] <= 16'h0430;
rommem[2321] <= 16'h3B43;
rommem[2322] <= 16'h0432;
rommem[2323] <= 16'h3B7C;
rommem[2324] <= 16'h0003;
rommem[2325] <= 16'h042E;
rommem[2326] <= 16'h5386;
rommem[2327] <= 16'h669E;
rommem[2328] <= 16'h4E75;
rommem[2329] <= 16'h4DF9;
rommem[2330] <= 16'hFFDC;
rommem[2331] <= 16'h0000;
rommem[2332] <= 16'h4BF9;
rommem[2333] <= 16'hFFE0;
rommem[2334] <= 16'h0000;
rommem[2335] <= 16'h2C3C;
rommem[2336] <= 16'h0003;
rommem[2337] <= 16'h0D40;
rommem[2338] <= 16'h33FC;
rommem[2339] <= 16'h000A;
rommem[2340] <= 16'hFFDC;
rommem[2341] <= 16'h0600;
rommem[2342] <= 16'h302D;
rommem[2343] <= 16'h04AC;
rommem[2344] <= 16'h0800;
rommem[2345] <= 16'h000E;
rommem[2346] <= 16'h6706;
rommem[2347] <= 16'h0800;
rommem[2348] <= 16'h000D;
rommem[2349] <= 16'h67E8;
rommem[2350] <= 16'h33FC;
rommem[2351] <= 16'h000B;
rommem[2352] <= 16'hFFDC;
rommem[2353] <= 16'h0600;
rommem[2354] <= 16'h202E;
rommem[2355] <= 16'h0C00;
rommem[2356] <= 16'h3200;
rommem[2357] <= 16'h4840;
rommem[2358] <= 16'h0240;
rommem[2359] <= 16'h00FF;
rommem[2360] <= 16'h0241;
rommem[2361] <= 16'h00FF;
rommem[2362] <= 16'h426E;
rommem[2363] <= 16'h0C04;
rommem[2364] <= 16'h242E;
rommem[2365] <= 16'h0C00;
rommem[2366] <= 16'h3602;
rommem[2367] <= 16'h4842;
rommem[2368] <= 16'h0242;
rommem[2369] <= 16'h00FF;
rommem[2370] <= 16'h0243;
rommem[2371] <= 16'h00FF;
rommem[2372] <= 16'h426E;
rommem[2373] <= 16'h0C04;
rommem[2374] <= 16'h282E;
rommem[2375] <= 16'h0C00;
rommem[2376] <= 16'h0244;
rommem[2377] <= 16'h7FFF;
rommem[2378] <= 16'h426E;
rommem[2379] <= 16'h0C04;
rommem[2380] <= 16'h3E2D;
rommem[2381] <= 16'h042C;
rommem[2382] <= 16'hBE7C;
rommem[2383] <= 16'h001C;
rommem[2384] <= 16'h64F6;
rommem[2385] <= 16'h33FC;
rommem[2386] <= 16'h000C;
rommem[2387] <= 16'hFFDC;
rommem[2388] <= 16'h0600;
rommem[2389] <= 16'h3B7C;
rommem[2390] <= 16'h0001;
rommem[2391] <= 16'h0422;
rommem[2392] <= 16'h3B44;
rommem[2393] <= 16'h0424;
rommem[2394] <= 16'h3B40;
rommem[2395] <= 16'h0426;
rommem[2396] <= 16'h3B41;
rommem[2397] <= 16'h0428;
rommem[2398] <= 16'h3B42;
rommem[2399] <= 16'h0430;
rommem[2400] <= 16'h3B43;
rommem[2401] <= 16'h0432;
rommem[2402] <= 16'h3B7C;
rommem[2403] <= 16'h0002;
rommem[2404] <= 16'h042E;
rommem[2405] <= 16'h5386;
rommem[2406] <= 16'h6600;
rommem[2407] <= 16'hFF76;
rommem[2408] <= 16'h4E75;
rommem[2409] <= 16'h4BF9;
rommem[2410] <= 16'hFFE0;
rommem[2411] <= 16'h0000;
rommem[2412] <= 16'h302D;
rommem[2413] <= 16'h04AC;
rommem[2414] <= 16'h0800;
rommem[2415] <= 16'h000D;
rommem[2416] <= 16'h67F6;
rommem[2417] <= 16'h2B7C;
rommem[2418] <= 16'h0000;
rommem[2419] <= 16'h1F40;
rommem[2420] <= 16'h04BC;
rommem[2421] <= 16'h3B7C;
rommem[2422] <= 16'h7C00;
rommem[2423] <= 16'h04A8;
rommem[2424] <= 16'h2B7C;
rommem[2425] <= 16'h0000;
rommem[2426] <= 16'h0118;
rommem[2427] <= 16'h0498;
rommem[2428] <= 16'h2B7C;
rommem[2429] <= 16'h0000;
rommem[2430] <= 16'h0028;
rommem[2431] <= 16'h04A4;
rommem[2432] <= 16'h2B7C;
rommem[2433] <= 16'h0000;
rommem[2434] <= 16'h0118;
rommem[2435] <= 16'h049C;
rommem[2436] <= 16'h3B7C;
rommem[2437] <= 16'h8080;
rommem[2438] <= 16'h04AC;
rommem[2439] <= 16'h302D;
rommem[2440] <= 16'h04AC;
rommem[2441] <= 16'h0800;
rommem[2442] <= 16'h000D;
rommem[2443] <= 16'h67F6;
rommem[2444] <= 16'h2B7C;
rommem[2445] <= 16'h0000;
rommem[2446] <= 16'h03E8;
rommem[2447] <= 16'h04B0;
rommem[2448] <= 16'h2B7C;
rommem[2449] <= 16'h0000;
rommem[2450] <= 16'h0000;
rommem[2451] <= 16'h0480;
rommem[2452] <= 16'h2B7C;
rommem[2453] <= 16'h0000;
rommem[2454] <= 16'h0118;
rommem[2455] <= 16'h0484;
rommem[2456] <= 16'h2B7C;
rommem[2457] <= 16'h0000;
rommem[2458] <= 16'h03E8;
rommem[2459] <= 16'h04B8;
rommem[2460] <= 16'h2B7C;
rommem[2461] <= 16'h0000;
rommem[2462] <= 16'h0000;
rommem[2463] <= 16'h0490;
rommem[2464] <= 16'h2B7C;
rommem[2465] <= 16'h0000;
rommem[2466] <= 16'h0118;
rommem[2467] <= 16'h0494;
rommem[2468] <= 16'h2B7C;
rommem[2469] <= 16'h0000;
rommem[2470] <= 16'h1F40;
rommem[2471] <= 16'h04BC;
rommem[2472] <= 16'h2B7C;
rommem[2473] <= 16'h0000;
rommem[2474] <= 16'h00F0;
rommem[2475] <= 16'h0498;
rommem[2476] <= 16'h2B7C;
rommem[2477] <= 16'h0000;
rommem[2478] <= 16'h0118;
rommem[2479] <= 16'h049C;
rommem[2480] <= 16'h2B7C;
rommem[2481] <= 16'h0000;
rommem[2482] <= 16'h0028;
rommem[2483] <= 16'h04A0;
rommem[2484] <= 16'h2B7C;
rommem[2485] <= 16'h0000;
rommem[2486] <= 16'h0028;
rommem[2487] <= 16'h04A4;
rommem[2488] <= 16'h3B7C;
rommem[2489] <= 16'h0091;
rommem[2490] <= 16'h04AE;
rommem[2491] <= 16'h3B7C;
rommem[2492] <= 16'h80A2;
rommem[2493] <= 16'h04AC;
rommem[2494] <= 16'h302D;
rommem[2495] <= 16'h04AC;
rommem[2496] <= 16'h0800;
rommem[2497] <= 16'h000D;
rommem[2498] <= 16'h67F6;
rommem[2499] <= 16'h4E75;
rommem[2500] <= 16'h4DF9;
rommem[2501] <= 16'hFFDC;
rommem[2502] <= 16'h0E00;
rommem[2503] <= 16'h3CBC;
rommem[2504] <= 16'h0013;
rommem[2505] <= 16'h3D7C;
rommem[2506] <= 16'h0000;
rommem[2507] <= 16'h0002;
rommem[2508] <= 16'h4DF9;
rommem[2509] <= 16'hFFDC;
rommem[2510] <= 16'h0E10;
rommem[2511] <= 16'h3CBC;
rommem[2512] <= 16'h0013;
rommem[2513] <= 16'h3D7C;
rommem[2514] <= 16'h0000;
rommem[2515] <= 16'h0002;
rommem[2516] <= 16'h4E75;
rommem[2517] <= 16'h3F00;
rommem[2518] <= 16'h302E;
rommem[2519] <= 16'h000A;
rommem[2520] <= 16'h0800;
rommem[2521] <= 16'h0001;
rommem[2522] <= 16'h66F6;
rommem[2523] <= 16'h301F;
rommem[2524] <= 16'h4E75;
rommem[2525] <= 16'h3D40;
rommem[2526] <= 16'h0006;
rommem[2527] <= 16'h3D41;
rommem[2528] <= 16'h0008;
rommem[2529] <= 16'h6100;
rommem[2530] <= 16'hFFE6;
rommem[2531] <= 16'h302E;
rommem[2532] <= 16'h000A;
rommem[2533] <= 16'h4E75;
rommem[2534] <= 16'h3F00;
rommem[2535] <= 16'h3D7C;
rommem[2536] <= 16'h0001;
rommem[2537] <= 16'h0004;
rommem[2538] <= 16'h7076;
rommem[2539] <= 16'h323C;
rommem[2540] <= 16'h0090;
rommem[2541] <= 16'h6100;
rommem[2542] <= 16'hFFDE;
rommem[2543] <= 16'h6100;
rommem[2544] <= 16'h0010;
rommem[2545] <= 16'h301F;
rommem[2546] <= 16'h323C;
rommem[2547] <= 16'h0050;
rommem[2548] <= 16'h6100;
rommem[2549] <= 16'hFFD0;
rommem[2550] <= 16'h6100;
rommem[2551] <= 16'h0002;
rommem[2552] <= 16'h3F00;
rommem[2553] <= 16'h302E;
rommem[2554] <= 16'h000A;
rommem[2555] <= 16'h0800;
rommem[2556] <= 16'h0007;
rommem[2557] <= 16'h66F6;
rommem[2558] <= 16'h301F;
rommem[2559] <= 16'h4E75;
rommem[2560] <= 16'h7000;
rommem[2561] <= 16'h720E;
rommem[2562] <= 16'h6100;
rommem[2563] <= 16'h001C;
rommem[2564] <= 16'h7002;
rommem[2565] <= 16'h41F9;
rommem[2566] <= 16'hFFFC;
rommem[2567] <= 16'h147C;
rommem[2568] <= 16'h6100;
rommem[2569] <= 16'h0076;
rommem[2570] <= 16'h4E75;
rommem[2571] <= 16'h4E75;
rommem[2572] <= 16'h6100;
rommem[2573] <= 16'hFFE6;
rommem[2574] <= 16'h6100;
rommem[2575] <= 16'hFFF8;
rommem[2576] <= 16'h4E75;
rommem[2577] <= 16'h4DF9;
rommem[2578] <= 16'hFFDC;
rommem[2579] <= 16'h0E00;
rommem[2580] <= 16'h3D7C;
rommem[2581] <= 16'h0001;
rommem[2582] <= 16'h0004;
rommem[2583] <= 16'h3D7C;
rommem[2584] <= 16'h0076;
rommem[2585] <= 16'h0006;
rommem[2586] <= 16'h3D7C;
rommem[2587] <= 16'h0090;
rommem[2588] <= 16'h0008;
rommem[2589] <= 16'h6100;
rommem[2590] <= 16'hFF6E;
rommem[2591] <= 16'h6100;
rommem[2592] <= 16'hFFB0;
rommem[2593] <= 16'h3D7C;
rommem[2594] <= 16'h0040;
rommem[2595] <= 16'h0006;
rommem[2596] <= 16'h3D7C;
rommem[2597] <= 16'h0010;
rommem[2598] <= 16'h0008;
rommem[2599] <= 16'h6100;
rommem[2600] <= 16'hFF5A;
rommem[2601] <= 16'h6100;
rommem[2602] <= 16'hFF9C;
rommem[2603] <= 16'h3D40;
rommem[2604] <= 16'h0006;
rommem[2605] <= 16'h3D7C;
rommem[2606] <= 16'h0010;
rommem[2607] <= 16'h0008;
rommem[2608] <= 16'h6100;
rommem[2609] <= 16'hFF48;
rommem[2610] <= 16'h6100;
rommem[2611] <= 16'hFF8A;
rommem[2612] <= 16'h3D41;
rommem[2613] <= 16'h0006;
rommem[2614] <= 16'h3D7C;
rommem[2615] <= 16'h0050;
rommem[2616] <= 16'h0008;
rommem[2617] <= 16'h6100;
rommem[2618] <= 16'hFF36;
rommem[2619] <= 16'h6100;
rommem[2620] <= 16'hFF78;
rommem[2621] <= 16'h4E75;
rommem[2622] <= 16'h0000;
rommem[2623] <= 16'h007D;
rommem[2624] <= 16'h0000;
rommem[2625] <= 16'h000C;
rommem[2626] <= 16'h0020;
rommem[2627] <= 16'h0001;
rommem[2628] <= 16'h41F9;
rommem[2629] <= 16'hFFFC;
rommem[2630] <= 16'h147C;
rommem[2631] <= 16'h4DF9;
rommem[2632] <= 16'hFFDC;
rommem[2633] <= 16'h0E00;
rommem[2634] <= 16'h3D7C;
rommem[2635] <= 16'h0001;
rommem[2636] <= 16'h0004;
rommem[2637] <= 16'h3D7C;
rommem[2638] <= 16'h0076;
rommem[2639] <= 16'h0006;
rommem[2640] <= 16'h3D7C;
rommem[2641] <= 16'h0090;
rommem[2642] <= 16'h0008;
rommem[2643] <= 16'h6100;
rommem[2644] <= 16'hFF02;
rommem[2645] <= 16'h6100;
rommem[2646] <= 16'hFF44;
rommem[2647] <= 16'h3D7C;
rommem[2648] <= 16'h0040;
rommem[2649] <= 16'h0006;
rommem[2650] <= 16'h3D7C;
rommem[2651] <= 16'h0010;
rommem[2652] <= 16'h0008;
rommem[2653] <= 16'h6100;
rommem[2654] <= 16'hFEEE;
rommem[2655] <= 16'h6100;
rommem[2656] <= 16'hFF30;
rommem[2657] <= 16'h3D40;
rommem[2658] <= 16'h0006;
rommem[2659] <= 16'h3D7C;
rommem[2660] <= 16'h0010;
rommem[2661] <= 16'h0008;
rommem[2662] <= 16'h6100;
rommem[2663] <= 16'hFEDC;
rommem[2664] <= 16'h6100;
rommem[2665] <= 16'hFF1E;
rommem[2666] <= 16'h3D58;
rommem[2667] <= 16'h0006;
rommem[2668] <= 16'h3D7C;
rommem[2669] <= 16'h0010;
rommem[2670] <= 16'h0008;
rommem[2671] <= 16'h6100;
rommem[2672] <= 16'hFECA;
rommem[2673] <= 16'h6100;
rommem[2674] <= 16'hFF0C;
rommem[2675] <= 16'h3D58;
rommem[2676] <= 16'h0006;
rommem[2677] <= 16'h3D7C;
rommem[2678] <= 16'h0010;
rommem[2679] <= 16'h0008;
rommem[2680] <= 16'h6100;
rommem[2681] <= 16'hFEB8;
rommem[2682] <= 16'h6100;
rommem[2683] <= 16'hFEFA;
rommem[2684] <= 16'h3D58;
rommem[2685] <= 16'h0006;
rommem[2686] <= 16'h3D7C;
rommem[2687] <= 16'h0010;
rommem[2688] <= 16'h0008;
rommem[2689] <= 16'h6100;
rommem[2690] <= 16'hFEA6;
rommem[2691] <= 16'h6100;
rommem[2692] <= 16'hFEE8;
rommem[2693] <= 16'h3D58;
rommem[2694] <= 16'h0006;
rommem[2695] <= 16'h3D7C;
rommem[2696] <= 16'h0010;
rommem[2697] <= 16'h0008;
rommem[2698] <= 16'h6100;
rommem[2699] <= 16'hFE94;
rommem[2700] <= 16'h6100;
rommem[2701] <= 16'hFED6;
rommem[2702] <= 16'h3D58;
rommem[2703] <= 16'h0006;
rommem[2704] <= 16'h3D7C;
rommem[2705] <= 16'h0010;
rommem[2706] <= 16'h0008;
rommem[2707] <= 16'h6100;
rommem[2708] <= 16'hFE82;
rommem[2709] <= 16'h6100;
rommem[2710] <= 16'hFEC4;
rommem[2711] <= 16'h3D58;
rommem[2712] <= 16'h0006;
rommem[2713] <= 16'h3D7C;
rommem[2714] <= 16'h0050;
rommem[2715] <= 16'h0008;
rommem[2716] <= 16'h6100;
rommem[2717] <= 16'hFE70;
rommem[2718] <= 16'h6100;
rommem[2719] <= 16'hFEB2;
rommem[2720] <= 16'h4E75;
rommem[2721] <= 16'h7021;
rommem[2722] <= 16'h7200;
rommem[2723] <= 16'h6100;
rommem[2724] <= 16'hFEDA;
rommem[2725] <= 16'h7020;
rommem[2726] <= 16'h6100;
rommem[2727] <= 16'hFED4;
rommem[2728] <= 16'h7023;
rommem[2729] <= 16'h323C;
rommem[2730] <= 16'h00E7;
rommem[2731] <= 16'h6100;
rommem[2732] <= 16'hFECA;
rommem[2733] <= 16'h7024;
rommem[2734] <= 16'h323C;
rommem[2735] <= 16'h00E7;
rommem[2736] <= 16'h6100;
rommem[2737] <= 16'hFEC0;
rommem[2738] <= 16'h4E75;
rommem[2739] <= 16'h2C7C;
rommem[2740] <= 16'hFFDC;
rommem[2741] <= 16'h0E10;
rommem[2742] <= 16'h4BF9;
rommem[2743] <= 16'h0001;
rommem[2744] <= 16'h0600;
rommem[2745] <= 16'h3D7C;
rommem[2746] <= 16'h0080;
rommem[2747] <= 16'h0004;
rommem[2748] <= 16'h303C;
rommem[2749] <= 16'h00DE;
rommem[2750] <= 16'h323C;
rommem[2751] <= 16'h0090;
rommem[2752] <= 16'h6100;
rommem[2753] <= 16'hFE38;
rommem[2754] <= 16'h4A00;
rommem[2755] <= 16'h6B72;
rommem[2756] <= 16'h303C;
rommem[2757] <= 16'h0000;
rommem[2758] <= 16'h323C;
rommem[2759] <= 16'h0010;
rommem[2760] <= 16'h6100;
rommem[2761] <= 16'hFE28;
rommem[2762] <= 16'h4A00;
rommem[2763] <= 16'h6B62;
rommem[2764] <= 16'h303C;
rommem[2765] <= 16'h00DF;
rommem[2766] <= 16'h323C;
rommem[2767] <= 16'h0090;
rommem[2768] <= 16'h6100;
rommem[2769] <= 16'hFE18;
rommem[2770] <= 16'h4A00;
rommem[2771] <= 16'h6B52;
rommem[2772] <= 16'h343C;
rommem[2773] <= 16'h0020;
rommem[2774] <= 16'h3D7C;
rommem[2775] <= 16'h0020;
rommem[2776] <= 16'h0008;
rommem[2777] <= 16'h6100;
rommem[2778] <= 16'hFDF6;
rommem[2779] <= 16'h6100;
rommem[2780] <= 16'hFE38;
rommem[2781] <= 16'h302E;
rommem[2782] <= 16'h000A;
rommem[2783] <= 16'h4A00;
rommem[2784] <= 16'h6B38;
rommem[2785] <= 16'h302E;
rommem[2786] <= 16'h0006;
rommem[2787] <= 16'h1B80;
rommem[2788] <= 16'h2000;
rommem[2789] <= 16'h5242;
rommem[2790] <= 16'hB47C;
rommem[2791] <= 16'h005F;
rommem[2792] <= 16'h66DA;
rommem[2793] <= 16'h3D7C;
rommem[2794] <= 16'h0068;
rommem[2795] <= 16'h0008;
rommem[2796] <= 16'h6100;
rommem[2797] <= 16'hFDD0;
rommem[2798] <= 16'h6100;
rommem[2799] <= 16'hFE12;
rommem[2800] <= 16'h302E;
rommem[2801] <= 16'h000A;
rommem[2802] <= 16'h4A00;
rommem[2803] <= 16'h6B12;
rommem[2804] <= 16'h302E;
rommem[2805] <= 16'h0006;
rommem[2806] <= 16'h1B80;
rommem[2807] <= 16'h2000;
rommem[2808] <= 16'h3D7C;
rommem[2809] <= 16'h0000;
rommem[2810] <= 16'h0004;
rommem[2811] <= 16'h7000;
rommem[2812] <= 16'h4E75;
rommem[2813] <= 16'h3D7C;
rommem[2814] <= 16'h0000;
rommem[2815] <= 16'h0004;
rommem[2816] <= 16'h4E75;
rommem[2817] <= 16'h2C7C;
rommem[2818] <= 16'hFFDC;
rommem[2819] <= 16'h0E10;
rommem[2820] <= 16'h4BF9;
rommem[2821] <= 16'h0001;
rommem[2822] <= 16'h0600;
rommem[2823] <= 16'h3D7C;
rommem[2824] <= 16'h0080;
rommem[2825] <= 16'h0004;
rommem[2826] <= 16'h303C;
rommem[2827] <= 16'h00DE;
rommem[2828] <= 16'h323C;
rommem[2829] <= 16'h0090;
rommem[2830] <= 16'h6100;
rommem[2831] <= 16'hFD9C;
rommem[2832] <= 16'h4A00;
rommem[2833] <= 16'h6B46;
rommem[2834] <= 16'h303C;
rommem[2835] <= 16'h0000;
rommem[2836] <= 16'h323C;
rommem[2837] <= 16'h0010;
rommem[2838] <= 16'h6100;
rommem[2839] <= 16'hFD8C;
rommem[2840] <= 16'h4A00;
rommem[2841] <= 16'h6B36;
rommem[2842] <= 16'h343C;
rommem[2843] <= 16'h0020;
rommem[2844] <= 16'h1035;
rommem[2845] <= 16'h2000;
rommem[2846] <= 16'h323C;
rommem[2847] <= 16'h0010;
rommem[2848] <= 16'h6100;
rommem[2849] <= 16'hFD78;
rommem[2850] <= 16'h4A00;
rommem[2851] <= 16'h6B22;
rommem[2852] <= 16'h5242;
rommem[2853] <= 16'hB47C;
rommem[2854] <= 16'h005F;
rommem[2855] <= 16'h66E8;
rommem[2856] <= 16'h1035;
rommem[2857] <= 16'h2000;
rommem[2858] <= 16'h323C;
rommem[2859] <= 16'h0050;
rommem[2860] <= 16'h6100;
rommem[2861] <= 16'hFD60;
rommem[2862] <= 16'h4A00;
rommem[2863] <= 16'h6B0A;
rommem[2864] <= 16'h3D7C;
rommem[2865] <= 16'h0000;
rommem[2866] <= 16'h0004;
rommem[2867] <= 16'h7000;
rommem[2868] <= 16'h4E75;
rommem[2869] <= 16'h3D7C;
rommem[2870] <= 16'h0000;
rommem[2871] <= 16'h0004;
rommem[2872] <= 16'h4E75;
rommem[2873] <= 16'h5254;
rommem[2874] <= 16'h4320;
rommem[2875] <= 16'h7265;
rommem[2876] <= 16'h6164;
rommem[2877] <= 16'h2F77;
rommem[2878] <= 16'h7269;
rommem[2879] <= 16'h7465;
rommem[2880] <= 16'h2066;
rommem[2881] <= 16'h6169;
rommem[2882] <= 16'h6C65;
rommem[2883] <= 16'h642E;
rommem[2884] <= 16'h0D0A;
rommem[2885] <= 16'h004E;
rommem[2886] <= 16'h3456;
rommem[2887] <= 16'h2036;
rommem[2888] <= 16'h386B;
rommem[2889] <= 16'h2053;
rommem[2890] <= 16'h7973;
rommem[2891] <= 16'h7465;
rommem[2892] <= 16'h6D20;
rommem[2893] <= 16'h5374;
rommem[2894] <= 16'h6172;
rommem[2895] <= 16'h7469;
rommem[2896] <= 16'h6E67;
rommem[2897] <= 16'h0000;
rommem[2898] <= 16'h0000;
rommem[2899] <= 16'h0000;
rommem[2900] <= 16'h0000;
rommem[2901] <= 16'h0000;
rommem[2902] <= 16'h0000;
rommem[2903] <= 16'h0000;
rommem[2904] <= 16'h0000;
rommem[2905] <= 16'h0000;
rommem[2906] <= 16'h0000;
rommem[2907] <= 16'h0000;
rommem[2908] <= 16'h0000;
rommem[2909] <= 16'h0000;
rommem[2910] <= 16'h0000;
rommem[2911] <= 16'h0000;
rommem[2912] <= 16'h0000;
rommem[2913] <= 16'h0000;
rommem[2914] <= 16'h0000;
rommem[2915] <= 16'h0000;
rommem[2916] <= 16'h0000;
rommem[2917] <= 16'h0000;
rommem[2918] <= 16'h0000;
rommem[2919] <= 16'h0000;
rommem[2920] <= 16'h0000;
rommem[2921] <= 16'h0000;
rommem[2922] <= 16'h0000;
rommem[2923] <= 16'h0000;
rommem[2924] <= 16'h0000;
rommem[2925] <= 16'h0000;
rommem[2926] <= 16'h0000;
rommem[2927] <= 16'h0000;
rommem[2928] <= 16'h0000;
rommem[2929] <= 16'h0000;
rommem[2930] <= 16'h0000;
rommem[2931] <= 16'h0000;
rommem[2932] <= 16'h0000;
rommem[2933] <= 16'h0000;
rommem[2934] <= 16'h0000;
rommem[2935] <= 16'h0000;
rommem[2936] <= 16'h0000;
rommem[2937] <= 16'h0000;
rommem[2938] <= 16'h0000;
rommem[2939] <= 16'h0000;
rommem[2940] <= 16'h0000;
rommem[2941] <= 16'h0000;
rommem[2942] <= 16'h0000;
rommem[2943] <= 16'h0000;
rommem[2944] <= 16'h0000;
rommem[2945] <= 16'h0000;
rommem[2946] <= 16'h0000;
rommem[2947] <= 16'h0000;
rommem[2948] <= 16'h0000;
rommem[2949] <= 16'h0000;
rommem[2950] <= 16'h0000;
rommem[2951] <= 16'h0000;
rommem[2952] <= 16'h0000;
rommem[2953] <= 16'h0000;
rommem[2954] <= 16'h0000;
rommem[2955] <= 16'h0000;
rommem[2956] <= 16'h0000;
rommem[2957] <= 16'h0000;
rommem[2958] <= 16'h0000;
rommem[2959] <= 16'h0000;
rommem[2960] <= 16'h0000;
rommem[2961] <= 16'h0000;
rommem[2962] <= 16'h0000;
rommem[2963] <= 16'h0000;
rommem[2964] <= 16'h0000;
rommem[2965] <= 16'h0000;
rommem[2966] <= 16'h0000;
rommem[2967] <= 16'h0000;
rommem[2968] <= 16'h0000;
rommem[2969] <= 16'h0000;
rommem[2970] <= 16'h0000;
rommem[2971] <= 16'h0000;
rommem[2972] <= 16'h0000;
rommem[2973] <= 16'h0000;
rommem[2974] <= 16'h0000;
rommem[2975] <= 16'h0000;
rommem[2976] <= 16'h0000;
rommem[2977] <= 16'h0000;
rommem[2978] <= 16'h0000;
rommem[2979] <= 16'h0000;
rommem[2980] <= 16'h0000;
rommem[2981] <= 16'h0000;
rommem[2982] <= 16'h0000;
rommem[2983] <= 16'h0000;
rommem[2984] <= 16'h0000;
rommem[2985] <= 16'h0000;
rommem[2986] <= 16'h0000;
rommem[2987] <= 16'h0000;
rommem[2988] <= 16'h0000;
rommem[2989] <= 16'h0000;
rommem[2990] <= 16'h0000;
rommem[2991] <= 16'h0000;
rommem[2992] <= 16'h0000;
rommem[2993] <= 16'h0000;
rommem[2994] <= 16'h0000;
rommem[2995] <= 16'h0000;
rommem[2996] <= 16'h0000;
rommem[2997] <= 16'h0000;
rommem[2998] <= 16'h0000;
rommem[2999] <= 16'h0000;
rommem[3000] <= 16'h0000;
rommem[3001] <= 16'h0000;
rommem[3002] <= 16'h0000;
rommem[3003] <= 16'h0000;
rommem[3004] <= 16'h0000;
rommem[3005] <= 16'h0000;
rommem[3006] <= 16'h0000;
rommem[3007] <= 16'h0000;
rommem[3008] <= 16'h0000;
rommem[3009] <= 16'h0000;
rommem[3010] <= 16'h0000;
rommem[3011] <= 16'h0000;
rommem[3012] <= 16'h0000;
rommem[3013] <= 16'h0000;
rommem[3014] <= 16'h0000;
rommem[3015] <= 16'h0000;
rommem[3016] <= 16'h0000;
rommem[3017] <= 16'h0000;
rommem[3018] <= 16'h0000;
rommem[3019] <= 16'h0000;
rommem[3020] <= 16'h0000;
rommem[3021] <= 16'h0000;
rommem[3022] <= 16'h0000;
rommem[3023] <= 16'h0000;
rommem[3024] <= 16'h0000;
rommem[3025] <= 16'h0000;
rommem[3026] <= 16'h0000;
rommem[3027] <= 16'h0000;
rommem[3028] <= 16'h0000;
rommem[3029] <= 16'h0018;
rommem[3030] <= 16'h1818;
rommem[3031] <= 16'h1818;
rommem[3032] <= 16'h0018;
rommem[3033] <= 16'h006C;
rommem[3034] <= 16'h6C00;
rommem[3035] <= 16'h0000;
rommem[3036] <= 16'h0000;
rommem[3037] <= 16'h006C;
rommem[3038] <= 16'h6CFE;
rommem[3039] <= 16'h6CFE;
rommem[3040] <= 16'h6C6C;
rommem[3041] <= 16'h0018;
rommem[3042] <= 16'h3E60;
rommem[3043] <= 16'h3C06;
rommem[3044] <= 16'h7C18;
rommem[3045] <= 16'h0000;
rommem[3046] <= 16'h66AC;
rommem[3047] <= 16'hD836;
rommem[3048] <= 16'h6ACC;
rommem[3049] <= 16'h0038;
rommem[3050] <= 16'h6C68;
rommem[3051] <= 16'h76DC;
rommem[3052] <= 16'hCE7B;
rommem[3053] <= 16'h0018;
rommem[3054] <= 16'h1830;
rommem[3055] <= 16'h0000;
rommem[3056] <= 16'h0000;
rommem[3057] <= 16'h000C;
rommem[3058] <= 16'h1830;
rommem[3059] <= 16'h3030;
rommem[3060] <= 16'h180C;
rommem[3061] <= 16'h0030;
rommem[3062] <= 16'h180C;
rommem[3063] <= 16'h0C0C;
rommem[3064] <= 16'h1830;
rommem[3065] <= 16'h0000;
rommem[3066] <= 16'h663C;
rommem[3067] <= 16'hFF3C;
rommem[3068] <= 16'h6600;
rommem[3069] <= 16'h0000;
rommem[3070] <= 16'h1818;
rommem[3071] <= 16'h7E18;
rommem[3072] <= 16'h1800;
rommem[3073] <= 16'h0000;
rommem[3074] <= 16'h0000;
rommem[3075] <= 16'h0000;
rommem[3076] <= 16'h1818;
rommem[3077] <= 16'h3000;
rommem[3078] <= 16'h0000;
rommem[3079] <= 16'h7E00;
rommem[3080] <= 16'h0000;
rommem[3081] <= 16'h0000;
rommem[3082] <= 16'h0000;
rommem[3083] <= 16'h0000;
rommem[3084] <= 16'h1818;
rommem[3085] <= 16'h0003;
rommem[3086] <= 16'h060C;
rommem[3087] <= 16'h1830;
rommem[3088] <= 16'h60C0;
rommem[3089] <= 16'h003C;
rommem[3090] <= 16'h666E;
rommem[3091] <= 16'h7E76;
rommem[3092] <= 16'h663C;
rommem[3093] <= 16'h0018;
rommem[3094] <= 16'h3878;
rommem[3095] <= 16'h1818;
rommem[3096] <= 16'h1818;
rommem[3097] <= 16'h003C;
rommem[3098] <= 16'h6606;
rommem[3099] <= 16'h0C18;
rommem[3100] <= 16'h307E;
rommem[3101] <= 16'h003C;
rommem[3102] <= 16'h6606;
rommem[3103] <= 16'h1C06;
rommem[3104] <= 16'h663C;
rommem[3105] <= 16'h001C;
rommem[3106] <= 16'h3C6C;
rommem[3107] <= 16'hCCFE;
rommem[3108] <= 16'h0C0C;
rommem[3109] <= 16'h007E;
rommem[3110] <= 16'h607C;
rommem[3111] <= 16'h0606;
rommem[3112] <= 16'h663C;
rommem[3113] <= 16'h001C;
rommem[3114] <= 16'h3060;
rommem[3115] <= 16'h7C66;
rommem[3116] <= 16'h663C;
rommem[3117] <= 16'h007E;
rommem[3118] <= 16'h0606;
rommem[3119] <= 16'h0C18;
rommem[3120] <= 16'h1818;
rommem[3121] <= 16'h003C;
rommem[3122] <= 16'h6666;
rommem[3123] <= 16'h3C66;
rommem[3124] <= 16'h663C;
rommem[3125] <= 16'h003C;
rommem[3126] <= 16'h6666;
rommem[3127] <= 16'h3E06;
rommem[3128] <= 16'h0C38;
rommem[3129] <= 16'h0000;
rommem[3130] <= 16'h1818;
rommem[3131] <= 16'h0000;
rommem[3132] <= 16'h1818;
rommem[3133] <= 16'h0000;
rommem[3134] <= 16'h1818;
rommem[3135] <= 16'h0000;
rommem[3136] <= 16'h1818;
rommem[3137] <= 16'h3000;
rommem[3138] <= 16'h0618;
rommem[3139] <= 16'h6018;
rommem[3140] <= 16'h0600;
rommem[3141] <= 16'h0000;
rommem[3142] <= 16'h007E;
rommem[3143] <= 16'h007E;
rommem[3144] <= 16'h0000;
rommem[3145] <= 16'h0000;
rommem[3146] <= 16'h6018;
rommem[3147] <= 16'h0618;
rommem[3148] <= 16'h6000;
rommem[3149] <= 16'h003C;
rommem[3150] <= 16'h6606;
rommem[3151] <= 16'h0C18;
rommem[3152] <= 16'h0018;
rommem[3153] <= 16'h007C;
rommem[3154] <= 16'hC6DE;
rommem[3155] <= 16'hD6DE;
rommem[3156] <= 16'hC078;
rommem[3157] <= 16'h003C;
rommem[3158] <= 16'h6666;
rommem[3159] <= 16'h7E66;
rommem[3160] <= 16'h6666;
rommem[3161] <= 16'h007C;
rommem[3162] <= 16'h6666;
rommem[3163] <= 16'h7C66;
rommem[3164] <= 16'h667C;
rommem[3165] <= 16'h001E;
rommem[3166] <= 16'h3060;
rommem[3167] <= 16'h6060;
rommem[3168] <= 16'h301E;
rommem[3169] <= 16'h0078;
rommem[3170] <= 16'h6C66;
rommem[3171] <= 16'h6666;
rommem[3172] <= 16'h6C78;
rommem[3173] <= 16'h007E;
rommem[3174] <= 16'h6060;
rommem[3175] <= 16'h7860;
rommem[3176] <= 16'h607E;
rommem[3177] <= 16'h007E;
rommem[3178] <= 16'h6060;
rommem[3179] <= 16'h7860;
rommem[3180] <= 16'h6060;
rommem[3181] <= 16'h003C;
rommem[3182] <= 16'h6660;
rommem[3183] <= 16'h6E66;
rommem[3184] <= 16'h663E;
rommem[3185] <= 16'h0066;
rommem[3186] <= 16'h6666;
rommem[3187] <= 16'h7E66;
rommem[3188] <= 16'h6666;
rommem[3189] <= 16'h003C;
rommem[3190] <= 16'h1818;
rommem[3191] <= 16'h1818;
rommem[3192] <= 16'h183C;
rommem[3193] <= 16'h0006;
rommem[3194] <= 16'h0606;
rommem[3195] <= 16'h0606;
rommem[3196] <= 16'h663C;
rommem[3197] <= 16'h00C6;
rommem[3198] <= 16'hCCD8;
rommem[3199] <= 16'hF0D8;
rommem[3200] <= 16'hCCC6;
rommem[3201] <= 16'h0060;
rommem[3202] <= 16'h6060;
rommem[3203] <= 16'h6060;
rommem[3204] <= 16'h607E;
rommem[3205] <= 16'h00C6;
rommem[3206] <= 16'hEEFE;
rommem[3207] <= 16'hD6C6;
rommem[3208] <= 16'hC6C6;
rommem[3209] <= 16'h00C6;
rommem[3210] <= 16'hE6F6;
rommem[3211] <= 16'hDECE;
rommem[3212] <= 16'hC6C6;
rommem[3213] <= 16'h003C;
rommem[3214] <= 16'h6666;
rommem[3215] <= 16'h6666;
rommem[3216] <= 16'h663C;
rommem[3217] <= 16'h007C;
rommem[3218] <= 16'h6666;
rommem[3219] <= 16'h7C60;
rommem[3220] <= 16'h6060;
rommem[3221] <= 16'h0078;
rommem[3222] <= 16'hCCCC;
rommem[3223] <= 16'hCCCC;
rommem[3224] <= 16'hDC7E;
rommem[3225] <= 16'h007C;
rommem[3226] <= 16'h6666;
rommem[3227] <= 16'h7C6C;
rommem[3228] <= 16'h6666;
rommem[3229] <= 16'h003C;
rommem[3230] <= 16'h6670;
rommem[3231] <= 16'h3C0E;
rommem[3232] <= 16'h663C;
rommem[3233] <= 16'h007E;
rommem[3234] <= 16'h1818;
rommem[3235] <= 16'h1818;
rommem[3236] <= 16'h1818;
rommem[3237] <= 16'h0066;
rommem[3238] <= 16'h6666;
rommem[3239] <= 16'h6666;
rommem[3240] <= 16'h663C;
rommem[3241] <= 16'h0066;
rommem[3242] <= 16'h6666;
rommem[3243] <= 16'h663C;
rommem[3244] <= 16'h3C18;
rommem[3245] <= 16'h00C6;
rommem[3246] <= 16'hC6C6;
rommem[3247] <= 16'hD6FE;
rommem[3248] <= 16'hEEC6;
rommem[3249] <= 16'h00C3;
rommem[3250] <= 16'h663C;
rommem[3251] <= 16'h183C;
rommem[3252] <= 16'h66C3;
rommem[3253] <= 16'h00C3;
rommem[3254] <= 16'h663C;
rommem[3255] <= 16'h1818;
rommem[3256] <= 16'h1818;
rommem[3257] <= 16'h00FE;
rommem[3258] <= 16'h0C18;
rommem[3259] <= 16'h3060;
rommem[3260] <= 16'hC0FE;
rommem[3261] <= 16'h003C;
rommem[3262] <= 16'h3030;
rommem[3263] <= 16'h3030;
rommem[3264] <= 16'h303C;
rommem[3265] <= 16'h00C0;
rommem[3266] <= 16'h6030;
rommem[3267] <= 16'h180C;
rommem[3268] <= 16'h0603;
rommem[3269] <= 16'h003C;
rommem[3270] <= 16'h0C0C;
rommem[3271] <= 16'h0C0C;
rommem[3272] <= 16'h0C3C;
rommem[3273] <= 16'h0010;
rommem[3274] <= 16'h386C;
rommem[3275] <= 16'hC600;
rommem[3276] <= 16'h0000;
rommem[3277] <= 16'h0000;
rommem[3278] <= 16'h0000;
rommem[3279] <= 16'h0000;
rommem[3280] <= 16'h0000;
rommem[3281] <= 16'hFE18;
rommem[3282] <= 16'h180C;
rommem[3283] <= 16'h0000;
rommem[3284] <= 16'h0000;
rommem[3285] <= 16'h0000;
rommem[3286] <= 16'h003C;
rommem[3287] <= 16'h063E;
rommem[3288] <= 16'h663E;
rommem[3289] <= 16'h0060;
rommem[3290] <= 16'h607C;
rommem[3291] <= 16'h6666;
rommem[3292] <= 16'h667C;
rommem[3293] <= 16'h0000;
rommem[3294] <= 16'h003C;
rommem[3295] <= 16'h6060;
rommem[3296] <= 16'h603C;
rommem[3297] <= 16'h0006;
rommem[3298] <= 16'h063E;
rommem[3299] <= 16'h6666;
rommem[3300] <= 16'h663E;
rommem[3301] <= 16'h0000;
rommem[3302] <= 16'h003C;
rommem[3303] <= 16'h667E;
rommem[3304] <= 16'h603C;
rommem[3305] <= 16'h001C;
rommem[3306] <= 16'h307C;
rommem[3307] <= 16'h3030;
rommem[3308] <= 16'h3030;
rommem[3309] <= 16'h0000;
rommem[3310] <= 16'h003E;
rommem[3311] <= 16'h6666;
rommem[3312] <= 16'h3E06;
rommem[3313] <= 16'h3C60;
rommem[3314] <= 16'h607C;
rommem[3315] <= 16'h6666;
rommem[3316] <= 16'h6666;
rommem[3317] <= 16'h0018;
rommem[3318] <= 16'h0018;
rommem[3319] <= 16'h1818;
rommem[3320] <= 16'h180C;
rommem[3321] <= 16'h000C;
rommem[3322] <= 16'h000C;
rommem[3323] <= 16'h0C0C;
rommem[3324] <= 16'h0C0C;
rommem[3325] <= 16'h7860;
rommem[3326] <= 16'h6066;
rommem[3327] <= 16'h6C78;
rommem[3328] <= 16'h6C66;
rommem[3329] <= 16'h0018;
rommem[3330] <= 16'h1818;
rommem[3331] <= 16'h1818;
rommem[3332] <= 16'h180C;
rommem[3333] <= 16'h0000;
rommem[3334] <= 16'h00EC;
rommem[3335] <= 16'hFED6;
rommem[3336] <= 16'hC6C6;
rommem[3337] <= 16'h0000;
rommem[3338] <= 16'h007C;
rommem[3339] <= 16'h6666;
rommem[3340] <= 16'h6666;
rommem[3341] <= 16'h0000;
rommem[3342] <= 16'h003C;
rommem[3343] <= 16'h6666;
rommem[3344] <= 16'h663C;
rommem[3345] <= 16'h0000;
rommem[3346] <= 16'h007C;
rommem[3347] <= 16'h6666;
rommem[3348] <= 16'h7C60;
rommem[3349] <= 16'h6000;
rommem[3350] <= 16'h003E;
rommem[3351] <= 16'h6666;
rommem[3352] <= 16'h3E06;
rommem[3353] <= 16'h0600;
rommem[3354] <= 16'h007C;
rommem[3355] <= 16'h6660;
rommem[3356] <= 16'h6060;
rommem[3357] <= 16'h0000;
rommem[3358] <= 16'h003C;
rommem[3359] <= 16'h603C;
rommem[3360] <= 16'h067C;
rommem[3361] <= 16'h0030;
rommem[3362] <= 16'h307C;
rommem[3363] <= 16'h3030;
rommem[3364] <= 16'h301C;
rommem[3365] <= 16'h0000;
rommem[3366] <= 16'h0066;
rommem[3367] <= 16'h6666;
rommem[3368] <= 16'h663E;
rommem[3369] <= 16'h0000;
rommem[3370] <= 16'h0066;
rommem[3371] <= 16'h6666;
rommem[3372] <= 16'h3C18;
rommem[3373] <= 16'h0000;
rommem[3374] <= 16'h00C6;
rommem[3375] <= 16'hC6D6;
rommem[3376] <= 16'hFE6C;
rommem[3377] <= 16'h0000;
rommem[3378] <= 16'h00C6;
rommem[3379] <= 16'h6C38;
rommem[3380] <= 16'h6CC6;
rommem[3381] <= 16'h0000;
rommem[3382] <= 16'h0066;
rommem[3383] <= 16'h6666;
rommem[3384] <= 16'h3C18;
rommem[3385] <= 16'h3000;
rommem[3386] <= 16'h007E;
rommem[3387] <= 16'h0C18;
rommem[3388] <= 16'h307E;
rommem[3389] <= 16'h000E;
rommem[3390] <= 16'h1818;
rommem[3391] <= 16'h7018;
rommem[3392] <= 16'h180E;
rommem[3393] <= 16'h0018;
rommem[3394] <= 16'h1818;
rommem[3395] <= 16'h1818;
rommem[3396] <= 16'h1818;
rommem[3397] <= 16'h0070;
rommem[3398] <= 16'h1818;
rommem[3399] <= 16'h0E18;
rommem[3400] <= 16'h1870;
rommem[3401] <= 16'h0072;
rommem[3402] <= 16'h9C00;
rommem[3403] <= 16'h0000;
rommem[3404] <= 16'h0000;
rommem[3405] <= 16'h00FE;
rommem[3406] <= 16'hFEFE;
rommem[3407] <= 16'hFEFE;
rommem[3408] <= 16'hFEFE;
