
module FT816_tb();

reg [5:0] btn;
reg clk;
always #10 clk <= ~clk;

initial begin
	#1 clk <= 1'b0;
	#50 btn <= 6'h00;
	#50 btn <= 6'h3F;
end

FT816Sys u1
(
	.btn(btn),
	.xclk(clk),
	.Led(),
	.sw(8'h00)
);

always @(posedge clk)
begin
	$display("%d %s", $time, u1.u1.u1.fnStateName(u1.u1.u1.state));
end

endmodule
