
module FT64_idissue();
endmodule
