`ifndef THOR2020_CONFIG_SV
`define THOR2020_CONFIG_SV

`define ABW		32
`define AMSB	31

`endif
