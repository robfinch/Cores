module redor32
(
	input [4:0] a,
	input [31:0] b,
	output reg o
);

	always @(a,b)
	case (a)
	5'd0:	o =  b[0];
	5'd1:	o = |b[1:0];
	5'd2:	o = |b[2:0];
	5'd3:	o = |b[3:0];
	5'd4:	o = |b[4:0];
	5'd5:	o = |b[5:0];
	5'd6:	o = |b[6:0];
	5'd7:	o = |b[7:0];
	5'd8:	o = |b[8:0];
	5'd9:	o = |b[9:0];
	5'd10:	o = |b[10:0];
	5'd11:	o = |b[11:0];
	5'd12:	o = |b[12:0];
	5'd13:	o = |b[13:0];
	5'd14:	o = |b[14:0];
	5'd15:	o = |b[15:0];
	5'd16:	o = |b[16:0];
	5'd17:	o = |b[17:0];
	5'd18:	o = |b[18:0];
	5'd19:	o = |b[19:0];
	5'd20:	o = |b[20:0];
	5'd21:	o = |b[21:0];
	5'd22:	o = |b[22:0];
	5'd23:	o = |b[23:0];
	5'd24:	o = |b[24:0];
	5'd25:	o = |b[25:0];
	5'd26:	o = |b[26:0];
	5'd27:	o = |b[27:0];
	5'd28:	o = |b[28:0];
	5'd29:	o = |b[29:0];
	5'd30:	o = |b[30:0];
	5'd31:	o = |b[31:0];
	endcase

endmodule
