`define AMSB  63
