parameter BIDLE = 5'd0;
parameter B_StoreAck = 5'd1;
parameter B_DCacheLoadStart = 5'd2;
parameter B_DCacheLoadStb = 5'd3;
parameter B_DCacheLoadWait1 = 5'd4;
parameter B_DCacheLoadWait2 = 5'd5;
parameter B_DCacheLoadResetBusy = 5'd6;
parameter B_ICacheAck = 5'd7;
parameter B8 = 5'd8;
parameter B_ICacheNack = 5'd9;
parameter B_ICacheNack2 = 5'd10;
parameter B11 = 5'd11;
parameter B12 = 5'd12;
parameter B_DLoadAck = 5'd13;
parameter B14 = 5'd14;
parameter B15 = 5'd15;
parameter B16 = 5'd16;
parameter B17 = 5'd17;
parameter B18 = 5'd18;
parameter B_LSNAck = 5'd19;
parameter B2a = 5'd20;
parameter B2b = 5'd21;
parameter B2c = 5'd22;
parameter B_DCacheLoadAck = 5'd23;
parameter B20 = 5'd24;
parameter B21 = 5'd25;
parameter B_DCacheLoadWait3 = 5'd26;
parameter B_LoadDesc = 5'd27;
parameter B_LoadDescStb = 5'd28;
parameter B_WaitSeg = 5'd29;
parameter B_DLoadNack = 5'd30;

parameter IDLE = 4'd0;
parameter IC1 = 4'd1;
parameter IC2 = 4'd2;
parameter IC3 = 4'd3;
parameter IC_WaitL2 = 4'd4;
parameter IC5 = 4'd5;
parameter IC6 = 4'd6;
parameter IC7 = 4'd7;
parameter IC_Next = 4'd8;
parameter IC9 = 4'd9;
parameter IC10 = 4'd10;
parameter IC3a = 4'd11;
