module redor128
(
	input [6:0] a,
	input [127:0] b,
	output reg o
);

	always @(a,b)
	case (a)
	7'd0:	o =  b[0];
	7'd1:	o = |b[1:0];
	7'd2:	o = |b[2:0];
	7'd3:	o = |b[3:0];
	7'd4:	o = |b[4:0];
	7'd5:	o = |b[5:0];
	7'd6:	o = |b[6:0];
	7'd7:	o = |b[7:0];
	7'd8:	o = |b[8:0];
	7'd9:	o = |b[9:0];
	7'd10:	o = |b[10:0];
	7'd11:	o = |b[11:0];
	7'd12:	o = |b[12:0];
	7'd13:	o = |b[13:0];
	7'd14:	o = |b[14:0];
	7'd15:	o = |b[15:0];
	7'd16:	o = |b[16:0];
	7'd17:	o = |b[17:0];
	7'd18:	o = |b[18:0];
	7'd19:	o = |b[19:0];
	7'd20:	o = |b[20:0];
	7'd21:	o = |b[21:0];
	7'd22:	o = |b[22:0];
	7'd23:	o = |b[23:0];
	7'd24:	o = |b[24:0];
	7'd25:	o = |b[25:0];
	7'd26:	o = |b[26:0];
	7'd27:	o = |b[27:0];
	7'd28:	o = |b[28:0];
	7'd29:	o = |b[29:0];
	7'd30:	o = |b[30:0];
	7'd31:	o = |b[31:0];
	7'd32:	o = |b[32:0];
	7'd33:	o = |b[33:0];
	7'd34:	o = |b[34:0];
	7'd35:	o = |b[35:0];
	7'd36:	o = |b[36:0];
	7'd37:	o = |b[37:0];
	7'd38:	o = |b[38:0];
	7'd39:	o = |b[39:0];
	7'd40:	o = |b[40:0];
	7'd41:	o = |b[41:0];
	7'd42:	o = |b[42:0];
	7'd43:	o = |b[43:0];
	7'd44:	o = |b[44:0];
	7'd45:	o = |b[45:0];
	7'd46:	o = |b[46:0];
	7'd47:	o = |b[47:0];
	7'd48:	o = |b[48:0];
	7'd49:	o = |b[49:0];
	7'd50:	o = |b[50:0];
	7'd51:	o = |b[51:0];
	7'd52:	o = |b[52:0];
	7'd53:	o = |b[53:0];
	7'd54:	o = |b[54:0];
	7'd55:	o = |b[55:0];
	7'd56:	o = |b[56:0];
	7'd57:	o = |b[57:0];
	7'd58:	o = |b[58:0];
	7'd59:	o = |b[59:0];
	7'd60:	o = |b[60:0];
	7'd61:	o = |b[61:0];
	7'd62:	o = |b[62:0];
	7'd63:	o = |b[63:0];
	
	7'd64:	o =  |b[64:0];
    7'd65:    o = |b[65:0];
    7'd66:    o = |b[66:0];
    7'd67:    o = |b[67:0];
    7'd68:    o = |b[68:0];
    7'd69:    o = |b[69:0];
    7'd70:    o = |b[70:0];
    7'd71:    o = |b[71:0];
    7'd72:    o = |b[72:0];
    7'd73:    o = |b[73:0];
    7'd74:    o = |b[74:0];
    7'd75:    o = |b[75:0];
    7'd76:    o = |b[76:0];
    7'd77:    o = |b[77:0];
    7'd78:    o = |b[78:0];
    7'd79:    o = |b[79:0];
    7'd80:    o = |b[80:0];
    7'd81:    o = |b[81:0];
    7'd82:    o = |b[82:0];
    7'd83:    o = |b[83:0];
    7'd84:    o = |b[84:0];
    7'd85:    o = |b[85:0];
    7'd86:    o = |b[86:0];
    7'd87:    o = |b[87:0];
    7'd88:    o = |b[88:0];
    7'd89:    o = |b[89:0];
    7'd90:    o = |b[90:0];
    7'd91:    o = |b[91:0];
    7'd92:    o = |b[92:0];
    7'd93:    o = |b[93:0];
    7'd94:    o = |b[94:0];
    7'd95:    o = |b[95:0];
    7'd96:    o = |b[96:0];
    7'd97:    o = |b[97:0];
    7'd98:    o = |b[98:0];
    7'd99:    o = |b[99:0];
    7'd100:    o = |b[100:0];
    7'd101:    o = |b[101:0];
    7'd102:    o = |b[102:0];
    7'd103:    o = |b[103:0];
    7'd104:    o = |b[104:0];
    7'd105:    o = |b[105:0];
    7'd106:    o = |b[106:0];
    7'd107:    o = |b[107:0];
    7'd108:    o = |b[108:0];
    7'd109:    o = |b[109:0];
    7'd110:    o = |b[110:0];
    7'd111:    o = |b[111:0];
    7'd112:    o = |b[112:0];
    7'd113:    o = |b[113:0];
    7'd114:    o = |b[114:0];
    7'd115:    o = |b[115:0];
    7'd116:    o = |b[116:0];
    7'd117:    o = |b[117:0];
    7'd118:    o = |b[118:0];
    7'd119:    o = |b[119:0];
    7'd120:    o = |b[120:0];
    7'd121:    o = |b[121:0];
    7'd122:    o = |b[122:0];
    7'd123:    o = |b[123:0];
    7'd124:    o = |b[124:0];
    7'd125:    o = |b[125:0];
    7'd126:    o = |b[126:0];
    7'd127:    o = |b[127:0];
	endcase

endmodule
