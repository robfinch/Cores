
typedef logic [FPWID-1:0] tPosit;
