rommem[0] <= 16'h0001;
rommem[1] <= 16'h0000;
rommem[2] <= 16'hFFFF;
rommem[3] <= 16'h0010;
rommem[4] <= 16'h4141;
rommem[5] <= 16'h3030;
rommem[6] <= 16'h3030;
rommem[7] <= 16'h3030;
rommem[8] <= 16'h33FC;
rommem[9] <= 16'hA1A1;
rommem[10] <= 16'hFFDC;
rommem[11] <= 16'h0600;
rommem[12] <= 16'h7000;
rommem[13] <= 16'h7200;
rommem[14] <= 16'h7400;
rommem[15] <= 16'h7600;
rommem[16] <= 16'h7800;
rommem[17] <= 16'h7A00;
rommem[18] <= 16'h7C00;
rommem[19] <= 16'h7E00;
rommem[20] <= 16'h4288;
rommem[21] <= 16'h4289;
rommem[22] <= 16'h428A;
rommem[23] <= 16'h428B;
rommem[24] <= 16'h428C;
rommem[25] <= 16'h428D;
rommem[26] <= 16'h428E;
rommem[27] <= 16'h4E67;
rommem[28] <= 16'h4DF9;
rommem[29] <= 16'hFFDC;
rommem[30] <= 16'h0000;
rommem[31] <= 16'h426E;
rommem[32] <= 16'h0C06;
rommem[33] <= 16'h2D7C;
rommem[34] <= 16'h8888;
rommem[35] <= 16'h8888;
rommem[36] <= 16'h0C08;
rommem[37] <= 16'h2D7C;
rommem[38] <= 16'h0123;
rommem[39] <= 16'h4567;
rommem[40] <= 16'h0C0C;
rommem[41] <= 16'h207C;
rommem[42] <= 16'hFF80;
rommem[43] <= 16'h0000;
rommem[44] <= 16'h203C;
rommem[45] <= 16'h0000;
rommem[46] <= 16'h00DF;
rommem[47] <= 16'h223C;
rommem[48] <= 16'h0005;
rommem[49] <= 16'h0000;
rommem[50] <= 16'h202E;
rommem[51] <= 16'h0C00;
rommem[52] <= 16'h426E;
rommem[53] <= 16'h0C04;
rommem[54] <= 16'h30C0;
rommem[55] <= 16'h5381;
rommem[56] <= 16'h66F2;
rommem[57] <= 16'h33FC;
rommem[58] <= 16'hA2A2;
rommem[59] <= 16'hFFDC;
rommem[60] <= 16'h0600;
rommem[61] <= 16'h41F9;
rommem[62] <= 16'hFFFF;
rommem[63] <= 16'h0254;
rommem[64] <= 16'h223C;
rommem[65] <= 16'h0000;
rommem[66] <= 16'h1000;
rommem[67] <= 16'h227C;
rommem[68] <= 16'hFF97;
rommem[69] <= 16'h0000;
rommem[70] <= 16'h247C;
rommem[71] <= 16'hFF80;
rommem[72] <= 16'h0000;
rommem[73] <= 16'h7000;
rommem[74] <= 16'h1018;
rommem[75] <= 16'h32C0;
rommem[76] <= 16'h51C9;
rommem[77] <= 16'hFFFA;
rommem[78] <= 16'h33FC;
rommem[79] <= 16'hA3A3;
rommem[80] <= 16'hFFDC;
rommem[81] <= 16'h0600;
rommem[82] <= 16'h41F9;
rommem[83] <= 16'hFFFF;
rommem[84] <= 16'h023C;
rommem[85] <= 16'h247C;
rommem[86] <= 16'h1FFF;
rommem[87] <= 16'h0000;
rommem[88] <= 16'h227C;
rommem[89] <= 16'hFFE0;
rommem[90] <= 16'h0000;
rommem[91] <= 16'h7200;
rommem[92] <= 16'h7400;
rommem[93] <= 16'h3029;
rommem[94] <= 16'h042A;
rommem[95] <= 16'hB07C;
rommem[96] <= 16'h001C;
rommem[97] <= 16'h64F6;
rommem[98] <= 16'h1018;
rommem[99] <= 16'h6726;
rommem[100] <= 16'h48C0;
rommem[101] <= 16'h14C0;
rommem[102] <= 16'h3340;
rommem[103] <= 16'h0420;
rommem[104] <= 16'h337C;
rommem[105] <= 16'h01FF;
rommem[106] <= 16'h0422;
rommem[107] <= 16'h337C;
rommem[108] <= 16'h0003;
rommem[109] <= 16'h0424;
rommem[110] <= 16'h3341;
rommem[111] <= 16'h0426;
rommem[112] <= 16'h3342;
rommem[113] <= 16'h0428;
rommem[114] <= 16'h337C;
rommem[115] <= 16'h0000;
rommem[116] <= 16'h042E;
rommem[117] <= 16'h5041;
rommem[118] <= 16'h60CC;
rommem[119] <= 16'h33FC;
rommem[120] <= 16'hA4A4;
rommem[121] <= 16'hFFDC;
rommem[122] <= 16'h0600;
rommem[123] <= 16'h47F9;
rommem[124] <= 16'hFFFF;
rommem[125] <= 16'h00FE;
rommem[126] <= 16'h605E;
rommem[127] <= 16'h60FE;
rommem[128] <= 16'h33FC;
rommem[129] <= 16'hA6A6;
rommem[130] <= 16'hFFDC;
rommem[131] <= 16'h0600;
rommem[132] <= 16'h2C7C;
rommem[133] <= 16'hFFE0;
rommem[134] <= 16'h0000;
rommem[135] <= 16'h343C;
rommem[136] <= 16'h0007;
rommem[137] <= 16'h1001;
rommem[138] <= 16'h0240;
rommem[139] <= 16'h000F;
rommem[140] <= 16'h0C40;
rommem[141] <= 16'h0009;
rommem[142] <= 16'h6302;
rommem[143] <= 16'h5E40;
rommem[144] <= 16'h0640;
rommem[145] <= 16'h0030;
rommem[146] <= 16'h3602;
rommem[147] <= 16'hE743;
rommem[148] <= 16'h382E;
rommem[149] <= 16'h042A;
rommem[150] <= 16'hB87C;
rommem[151] <= 16'h001C;
rommem[152] <= 16'h64F6;
rommem[153] <= 16'h48C0;
rommem[154] <= 16'h3D40;
rommem[155] <= 16'h0420;
rommem[156] <= 16'h3D7C;
rommem[157] <= 16'h01FF;
rommem[158] <= 16'h0422;
rommem[159] <= 16'h3D7C;
rommem[160] <= 16'h0003;
rommem[161] <= 16'h0424;
rommem[162] <= 16'h3D43;
rommem[163] <= 16'h0426;
rommem[164] <= 16'h3D7C;
rommem[165] <= 16'h0008;
rommem[166] <= 16'h0428;
rommem[167] <= 16'h3D7C;
rommem[168] <= 16'h0000;
rommem[169] <= 16'h042E;
rommem[170] <= 16'hE899;
rommem[171] <= 16'h57CA;
rommem[172] <= 16'hFFBA;
rommem[173] <= 16'h4ED5;
rommem[174] <= 16'h33FC;
rommem[175] <= 16'hA5A5;
rommem[176] <= 16'hFFDC;
rommem[177] <= 16'h0600;
rommem[178] <= 16'h207C;
rommem[179] <= 16'h0000;
rommem[180] <= 16'h0008;
rommem[181] <= 16'h203C;
rommem[182] <= 16'hAAAA;
rommem[183] <= 16'h5555;
rommem[184] <= 16'h20C0;
rommem[185] <= 16'h2208;
rommem[186] <= 16'h4A41;
rommem[187] <= 16'h6608;
rommem[188] <= 16'h4BF9;
rommem[189] <= 16'hFFFF;
rommem[190] <= 16'h0180;
rommem[191] <= 16'h6080;
rommem[192] <= 16'h33FC;
rommem[193] <= 16'hA9A9;
rommem[194] <= 16'hFFDC;
rommem[195] <= 16'h0600;
rommem[196] <= 16'hB1FC;
rommem[197] <= 16'h1FFF;
rommem[198] <= 16'hFFFC;
rommem[199] <= 16'h66E0;
rommem[200] <= 16'h33FC;
rommem[201] <= 16'hA7A7;
rommem[202] <= 16'hFFDC;
rommem[203] <= 16'h0600;
rommem[204] <= 16'h2448;
rommem[205] <= 16'h207C;
rommem[206] <= 16'h0000;
rommem[207] <= 16'h0008;
rommem[208] <= 16'h2018;
rommem[209] <= 16'hB5C8;
rommem[210] <= 16'h671A;
rommem[211] <= 16'h2208;
rommem[212] <= 16'h4A41;
rommem[213] <= 16'h660A;
rommem[214] <= 16'h4BF9;
rommem[215] <= 16'hFFFF;
rommem[216] <= 16'h01B6;
rommem[217] <= 16'h6000;
rommem[218] <= 16'hFF4C;
rommem[219] <= 16'h0C80;
rommem[220] <= 16'hAAAA;
rommem[221] <= 16'h5555;
rommem[222] <= 16'h67E2;
rommem[223] <= 16'h6678;
rommem[224] <= 16'h33FC;
rommem[225] <= 16'hA8A8;
rommem[226] <= 16'hFFDC;
rommem[227] <= 16'h0600;
rommem[228] <= 16'h207C;
rommem[229] <= 16'h0000;
rommem[230] <= 16'h0008;
rommem[231] <= 16'h203C;
rommem[232] <= 16'h5555;
rommem[233] <= 16'hAAAA;
rommem[234] <= 16'h20C0;
rommem[235] <= 16'h2208;
rommem[236] <= 16'h4A41;
rommem[237] <= 16'h660A;
rommem[238] <= 16'h4BF9;
rommem[239] <= 16'hFFFF;
rommem[240] <= 16'h01E6;
rommem[241] <= 16'h6000;
rommem[242] <= 16'hFF1C;
rommem[243] <= 16'hB1FC;
rommem[244] <= 16'h1FFF;
rommem[245] <= 16'hFFFC;
rommem[246] <= 16'h66E6;
rommem[247] <= 16'h2448;
rommem[248] <= 16'h207C;
rommem[249] <= 16'h0000;
rommem[250] <= 16'h0008;
rommem[251] <= 16'h2018;
rommem[252] <= 16'hB5C8;
rommem[253] <= 16'h671A;
rommem[254] <= 16'h2208;
rommem[255] <= 16'h4A41;
rommem[256] <= 16'h660A;
rommem[257] <= 16'h4BF9;
rommem[258] <= 16'h0000;
rommem[259] <= 16'h0000;
rommem[260] <= 16'h6000;
rommem[261] <= 16'hFEF6;
rommem[262] <= 16'h0C80;
rommem[263] <= 16'h5555;
rommem[264] <= 16'hAAAA;
rommem[265] <= 16'h67E2;
rommem[266] <= 16'h6622;
rommem[267] <= 16'h23C8;
rommem[268] <= 16'h0000;
rommem[269] <= 16'h0000;
rommem[270] <= 16'h91FC;
rommem[271] <= 16'h0000;
rommem[272] <= 16'h000C;
rommem[273] <= 16'h21C8;
rommem[274] <= 16'h0404;
rommem[275] <= 16'h21FC;
rommem[276] <= 16'h4652;
rommem[277] <= 16'h4545;
rommem[278] <= 16'h0400;
rommem[279] <= 16'h21FC;
rommem[280] <= 16'h0000;
rommem[281] <= 16'h0408;
rommem[282] <= 16'h0408;
rommem[283] <= 16'h4ED3;
rommem[284] <= 16'h4ED3;
rommem[285] <= 16'h60FC;
rommem[286] <= 16'h4E34;
rommem[287] <= 16'h5620;
rommem[288] <= 16'h3638;
rommem[289] <= 16'h6B20;
rommem[290] <= 16'h5379;
rommem[291] <= 16'h7374;
rommem[292] <= 16'h656D;
rommem[293] <= 16'h2053;
rommem[294] <= 16'h7461;
rommem[295] <= 16'h7274;
rommem[296] <= 16'h696E;
rommem[297] <= 16'h6700;
rommem[298] <= 16'h0000;
rommem[299] <= 16'h0000;
rommem[300] <= 16'h0000;
rommem[301] <= 16'h0000;
rommem[302] <= 16'h0000;
rommem[303] <= 16'h0000;
rommem[304] <= 16'h0000;
rommem[305] <= 16'h0000;
rommem[306] <= 16'h0000;
rommem[307] <= 16'h0000;
rommem[308] <= 16'h0000;
rommem[309] <= 16'h0000;
rommem[310] <= 16'h0000;
rommem[311] <= 16'h0000;
rommem[312] <= 16'h0000;
rommem[313] <= 16'h0000;
rommem[314] <= 16'h0000;
rommem[315] <= 16'h0000;
rommem[316] <= 16'h0000;
rommem[317] <= 16'h0000;
rommem[318] <= 16'h0000;
rommem[319] <= 16'h0000;
rommem[320] <= 16'h0000;
rommem[321] <= 16'h0000;
rommem[322] <= 16'h0000;
rommem[323] <= 16'h0000;
rommem[324] <= 16'h0000;
rommem[325] <= 16'h0000;
rommem[326] <= 16'h0000;
rommem[327] <= 16'h0000;
rommem[328] <= 16'h0000;
rommem[329] <= 16'h0000;
rommem[330] <= 16'h0000;
rommem[331] <= 16'h0000;
rommem[332] <= 16'h0000;
rommem[333] <= 16'h0000;
rommem[334] <= 16'h0000;
rommem[335] <= 16'h0000;
rommem[336] <= 16'h0000;
rommem[337] <= 16'h0000;
rommem[338] <= 16'h0000;
rommem[339] <= 16'h0000;
rommem[340] <= 16'h0000;
rommem[341] <= 16'h0000;
rommem[342] <= 16'h0000;
rommem[343] <= 16'h0000;
rommem[344] <= 16'h0000;
rommem[345] <= 16'h0000;
rommem[346] <= 16'h0000;
rommem[347] <= 16'h0000;
rommem[348] <= 16'h0000;
rommem[349] <= 16'h0000;
rommem[350] <= 16'h0000;
rommem[351] <= 16'h0000;
rommem[352] <= 16'h0000;
rommem[353] <= 16'h0000;
rommem[354] <= 16'h0000;
rommem[355] <= 16'h0000;
rommem[356] <= 16'h0000;
rommem[357] <= 16'h0000;
rommem[358] <= 16'h0000;
rommem[359] <= 16'h0000;
rommem[360] <= 16'h0000;
rommem[361] <= 16'h0000;
rommem[362] <= 16'h0000;
rommem[363] <= 16'h0000;
rommem[364] <= 16'h0000;
rommem[365] <= 16'h0000;
rommem[366] <= 16'h0000;
rommem[367] <= 16'h0000;
rommem[368] <= 16'h0000;
rommem[369] <= 16'h0000;
rommem[370] <= 16'h0000;
rommem[371] <= 16'h0000;
rommem[372] <= 16'h0000;
rommem[373] <= 16'h0000;
rommem[374] <= 16'h0000;
rommem[375] <= 16'h0000;
rommem[376] <= 16'h0000;
rommem[377] <= 16'h0000;
rommem[378] <= 16'h0000;
rommem[379] <= 16'h0000;
rommem[380] <= 16'h0000;
rommem[381] <= 16'h0000;
rommem[382] <= 16'h0000;
rommem[383] <= 16'h0000;
rommem[384] <= 16'h0000;
rommem[385] <= 16'h0000;
rommem[386] <= 16'h0000;
rommem[387] <= 16'h0000;
rommem[388] <= 16'h0000;
rommem[389] <= 16'h0000;
rommem[390] <= 16'h0000;
rommem[391] <= 16'h0000;
rommem[392] <= 16'h0000;
rommem[393] <= 16'h0000;
rommem[394] <= 16'h0000;
rommem[395] <= 16'h0000;
rommem[396] <= 16'h0000;
rommem[397] <= 16'h0000;
rommem[398] <= 16'h0000;
rommem[399] <= 16'h0000;
rommem[400] <= 16'h0000;
rommem[401] <= 16'h0000;
rommem[402] <= 16'h0000;
rommem[403] <= 16'h0000;
rommem[404] <= 16'h0000;
rommem[405] <= 16'h0000;
rommem[406] <= 16'h0000;
rommem[407] <= 16'h0000;
rommem[408] <= 16'h0000;
rommem[409] <= 16'h0000;
rommem[410] <= 16'h0000;
rommem[411] <= 16'h0000;
rommem[412] <= 16'h0000;
rommem[413] <= 16'h0000;
rommem[414] <= 16'h0000;
rommem[415] <= 16'h0000;
rommem[416] <= 16'h0000;
rommem[417] <= 16'h0000;
rommem[418] <= 16'h0000;
rommem[419] <= 16'h0000;
rommem[420] <= 16'h0000;
rommem[421] <= 16'h0000;
rommem[422] <= 16'h0000;
rommem[423] <= 16'h0000;
rommem[424] <= 16'h0000;
rommem[425] <= 16'h0000;
rommem[426] <= 16'h0000;
rommem[427] <= 16'h0000;
rommem[428] <= 16'h0000;
rommem[429] <= 16'h0000;
rommem[430] <= 16'h1818;
rommem[431] <= 16'h1818;
rommem[432] <= 16'h1800;
rommem[433] <= 16'h1800;
rommem[434] <= 16'h6C6C;
rommem[435] <= 16'h0000;
rommem[436] <= 16'h0000;
rommem[437] <= 16'h0000;
rommem[438] <= 16'h6C6C;
rommem[439] <= 16'hFE6C;
rommem[440] <= 16'hFE6C;
rommem[441] <= 16'h6C00;
rommem[442] <= 16'h183E;
rommem[443] <= 16'h603C;
rommem[444] <= 16'h067C;
rommem[445] <= 16'h1800;
rommem[446] <= 16'h0066;
rommem[447] <= 16'hACD8;
rommem[448] <= 16'h366A;
rommem[449] <= 16'hCC00;
rommem[450] <= 16'h386C;
rommem[451] <= 16'h6876;
rommem[452] <= 16'hDCCE;
rommem[453] <= 16'h7B00;
rommem[454] <= 16'h1818;
rommem[455] <= 16'h3000;
rommem[456] <= 16'h0000;
rommem[457] <= 16'h0000;
rommem[458] <= 16'h0C18;
rommem[459] <= 16'h3030;
rommem[460] <= 16'h3018;
rommem[461] <= 16'h0C00;
rommem[462] <= 16'h3018;
rommem[463] <= 16'h0C0C;
rommem[464] <= 16'h0C18;
rommem[465] <= 16'h3000;
rommem[466] <= 16'h0066;
rommem[467] <= 16'h3CFF;
rommem[468] <= 16'h3C66;
rommem[469] <= 16'h0000;
rommem[470] <= 16'h0018;
rommem[471] <= 16'h187E;
rommem[472] <= 16'h1818;
rommem[473] <= 16'h0000;
rommem[474] <= 16'h0000;
rommem[475] <= 16'h0000;
rommem[476] <= 16'h0018;
rommem[477] <= 16'h1830;
rommem[478] <= 16'h0000;
rommem[479] <= 16'h007E;
rommem[480] <= 16'h0000;
rommem[481] <= 16'h0000;
rommem[482] <= 16'h0000;
rommem[483] <= 16'h0000;
rommem[484] <= 16'h0018;
rommem[485] <= 16'h1800;
rommem[486] <= 16'h0306;
rommem[487] <= 16'h0C18;
rommem[488] <= 16'h3060;
rommem[489] <= 16'hC000;
rommem[490] <= 16'h3C66;
rommem[491] <= 16'h6E7E;
rommem[492] <= 16'h7666;
rommem[493] <= 16'h3C00;
rommem[494] <= 16'h1838;
rommem[495] <= 16'h7818;
rommem[496] <= 16'h1818;
rommem[497] <= 16'h1800;
rommem[498] <= 16'h3C66;
rommem[499] <= 16'h060C;
rommem[500] <= 16'h1830;
rommem[501] <= 16'h7E00;
rommem[502] <= 16'h3C66;
rommem[503] <= 16'h061C;
rommem[504] <= 16'h0666;
rommem[505] <= 16'h3C00;
rommem[506] <= 16'h1C3C;
rommem[507] <= 16'h6CCC;
rommem[508] <= 16'hFE0C;
rommem[509] <= 16'h0C00;
rommem[510] <= 16'h7E60;
rommem[511] <= 16'h7C06;
rommem[512] <= 16'h0666;
rommem[513] <= 16'h3C00;
rommem[514] <= 16'h1C30;
rommem[515] <= 16'h607C;
rommem[516] <= 16'h6666;
rommem[517] <= 16'h3C00;
rommem[518] <= 16'h7E06;
rommem[519] <= 16'h060C;
rommem[520] <= 16'h1818;
rommem[521] <= 16'h1800;
rommem[522] <= 16'h3C66;
rommem[523] <= 16'h663C;
rommem[524] <= 16'h6666;
rommem[525] <= 16'h3C00;
rommem[526] <= 16'h3C66;
rommem[527] <= 16'h663E;
rommem[528] <= 16'h060C;
rommem[529] <= 16'h3800;
rommem[530] <= 16'h0018;
rommem[531] <= 16'h1800;
rommem[532] <= 16'h0018;
rommem[533] <= 16'h1800;
rommem[534] <= 16'h0018;
rommem[535] <= 16'h1800;
rommem[536] <= 16'h0018;
rommem[537] <= 16'h1830;
rommem[538] <= 16'h0006;
rommem[539] <= 16'h1860;
rommem[540] <= 16'h1806;
rommem[541] <= 16'h0000;
rommem[542] <= 16'h0000;
rommem[543] <= 16'h7E00;
rommem[544] <= 16'h7E00;
rommem[545] <= 16'h0000;
rommem[546] <= 16'h0060;
rommem[547] <= 16'h1806;
rommem[548] <= 16'h1860;
rommem[549] <= 16'h0000;
rommem[550] <= 16'h3C66;
rommem[551] <= 16'h060C;
rommem[552] <= 16'h1800;
rommem[553] <= 16'h1800;
rommem[554] <= 16'h7CC6;
rommem[555] <= 16'hDED6;
rommem[556] <= 16'hDEC0;
rommem[557] <= 16'h7800;
rommem[558] <= 16'h3C66;
rommem[559] <= 16'h667E;
rommem[560] <= 16'h6666;
rommem[561] <= 16'h6600;
rommem[562] <= 16'h7C66;
rommem[563] <= 16'h667C;
rommem[564] <= 16'h6666;
rommem[565] <= 16'h7C00;
rommem[566] <= 16'h1E30;
rommem[567] <= 16'h6060;
rommem[568] <= 16'h6030;
rommem[569] <= 16'h1E00;
rommem[570] <= 16'h786C;
rommem[571] <= 16'h6666;
rommem[572] <= 16'h666C;
rommem[573] <= 16'h7800;
rommem[574] <= 16'h7E60;
rommem[575] <= 16'h6078;
rommem[576] <= 16'h6060;
rommem[577] <= 16'h7E00;
rommem[578] <= 16'h7E60;
rommem[579] <= 16'h6078;
rommem[580] <= 16'h6060;
rommem[581] <= 16'h6000;
rommem[582] <= 16'h3C66;
rommem[583] <= 16'h606E;
rommem[584] <= 16'h6666;
rommem[585] <= 16'h3E00;
rommem[586] <= 16'h6666;
rommem[587] <= 16'h667E;
rommem[588] <= 16'h6666;
rommem[589] <= 16'h6600;
rommem[590] <= 16'h3C18;
rommem[591] <= 16'h1818;
rommem[592] <= 16'h1818;
rommem[593] <= 16'h3C00;
rommem[594] <= 16'h0606;
rommem[595] <= 16'h0606;
rommem[596] <= 16'h0666;
rommem[597] <= 16'h3C00;
rommem[598] <= 16'hC6CC;
rommem[599] <= 16'hD8F0;
rommem[600] <= 16'hD8CC;
rommem[601] <= 16'hC600;
rommem[602] <= 16'h6060;
rommem[603] <= 16'h6060;
rommem[604] <= 16'h6060;
rommem[605] <= 16'h7E00;
rommem[606] <= 16'hC6EE;
rommem[607] <= 16'hFED6;
rommem[608] <= 16'hC6C6;
rommem[609] <= 16'hC600;
rommem[610] <= 16'hC6E6;
rommem[611] <= 16'hF6DE;
rommem[612] <= 16'hCEC6;
rommem[613] <= 16'hC600;
rommem[614] <= 16'h3C66;
rommem[615] <= 16'h6666;
rommem[616] <= 16'h6666;
rommem[617] <= 16'h3C00;
rommem[618] <= 16'h7C66;
rommem[619] <= 16'h667C;
rommem[620] <= 16'h6060;
rommem[621] <= 16'h6000;
rommem[622] <= 16'h78CC;
rommem[623] <= 16'hCCCC;
rommem[624] <= 16'hCCDC;
rommem[625] <= 16'h7E00;
rommem[626] <= 16'h7C66;
rommem[627] <= 16'h667C;
rommem[628] <= 16'h6C66;
rommem[629] <= 16'h6600;
rommem[630] <= 16'h3C66;
rommem[631] <= 16'h703C;
rommem[632] <= 16'h0E66;
rommem[633] <= 16'h3C00;
rommem[634] <= 16'h7E18;
rommem[635] <= 16'h1818;
rommem[636] <= 16'h1818;
rommem[637] <= 16'h1800;
rommem[638] <= 16'h6666;
rommem[639] <= 16'h6666;
rommem[640] <= 16'h6666;
rommem[641] <= 16'h3C00;
rommem[642] <= 16'h6666;
rommem[643] <= 16'h6666;
rommem[644] <= 16'h3C3C;
rommem[645] <= 16'h1800;
rommem[646] <= 16'hC6C6;
rommem[647] <= 16'hC6D6;
rommem[648] <= 16'hFEEE;
rommem[649] <= 16'hC600;
rommem[650] <= 16'hC366;
rommem[651] <= 16'h3C18;
rommem[652] <= 16'h3C66;
rommem[653] <= 16'hC300;
rommem[654] <= 16'hC366;
rommem[655] <= 16'h3C18;
rommem[656] <= 16'h1818;
rommem[657] <= 16'h1800;
rommem[658] <= 16'hFE0C;
rommem[659] <= 16'h1830;
rommem[660] <= 16'h60C0;
rommem[661] <= 16'hFE00;
rommem[662] <= 16'h3C30;
rommem[663] <= 16'h3030;
rommem[664] <= 16'h3030;
rommem[665] <= 16'h3C00;
rommem[666] <= 16'hC060;
rommem[667] <= 16'h3018;
rommem[668] <= 16'h0C06;
rommem[669] <= 16'h0300;
rommem[670] <= 16'h3C0C;
rommem[671] <= 16'h0C0C;
rommem[672] <= 16'h0C0C;
rommem[673] <= 16'h3C00;
rommem[674] <= 16'h1038;
rommem[675] <= 16'h6CC6;
rommem[676] <= 16'h0000;
rommem[677] <= 16'h0000;
rommem[678] <= 16'h0000;
rommem[679] <= 16'h0000;
rommem[680] <= 16'h0000;
rommem[681] <= 16'h00FE;
rommem[682] <= 16'h1818;
rommem[683] <= 16'h0C00;
rommem[684] <= 16'h0000;
rommem[685] <= 16'h0000;
rommem[686] <= 16'h0000;
rommem[687] <= 16'h3C06;
rommem[688] <= 16'h3E66;
rommem[689] <= 16'h3E00;
rommem[690] <= 16'h6060;
rommem[691] <= 16'h7C66;
rommem[692] <= 16'h6666;
rommem[693] <= 16'h7C00;
rommem[694] <= 16'h0000;
rommem[695] <= 16'h3C60;
rommem[696] <= 16'h6060;
rommem[697] <= 16'h3C00;
rommem[698] <= 16'h0606;
rommem[699] <= 16'h3E66;
rommem[700] <= 16'h6666;
rommem[701] <= 16'h3E00;
rommem[702] <= 16'h0000;
rommem[703] <= 16'h3C66;
rommem[704] <= 16'h7E60;
rommem[705] <= 16'h3C00;
rommem[706] <= 16'h1C30;
rommem[707] <= 16'h7C30;
rommem[708] <= 16'h3030;
rommem[709] <= 16'h3000;
rommem[710] <= 16'h0000;
rommem[711] <= 16'h3E66;
rommem[712] <= 16'h663E;
rommem[713] <= 16'h063C;
rommem[714] <= 16'h6060;
rommem[715] <= 16'h7C66;
rommem[716] <= 16'h6666;
rommem[717] <= 16'h6600;
rommem[718] <= 16'h1800;
rommem[719] <= 16'h1818;
rommem[720] <= 16'h1818;
rommem[721] <= 16'h0C00;
rommem[722] <= 16'h0C00;
rommem[723] <= 16'h0C0C;
rommem[724] <= 16'h0C0C;
rommem[725] <= 16'h0C78;
rommem[726] <= 16'h6060;
rommem[727] <= 16'h666C;
rommem[728] <= 16'h786C;
rommem[729] <= 16'h6600;
rommem[730] <= 16'h1818;
rommem[731] <= 16'h1818;
rommem[732] <= 16'h1818;
rommem[733] <= 16'h0C00;
rommem[734] <= 16'h0000;
rommem[735] <= 16'hECFE;
rommem[736] <= 16'hD6C6;
rommem[737] <= 16'hC600;
rommem[738] <= 16'h0000;
rommem[739] <= 16'h7C66;
rommem[740] <= 16'h6666;
rommem[741] <= 16'h6600;
rommem[742] <= 16'h0000;
rommem[743] <= 16'h3C66;
rommem[744] <= 16'h6666;
rommem[745] <= 16'h3C00;
rommem[746] <= 16'h0000;
rommem[747] <= 16'h7C66;
rommem[748] <= 16'h667C;
rommem[749] <= 16'h6060;
rommem[750] <= 16'h0000;
rommem[751] <= 16'h3E66;
rommem[752] <= 16'h663E;
rommem[753] <= 16'h0606;
rommem[754] <= 16'h0000;
rommem[755] <= 16'h7C66;
rommem[756] <= 16'h6060;
rommem[757] <= 16'h6000;
rommem[758] <= 16'h0000;
rommem[759] <= 16'h3C60;
rommem[760] <= 16'h3C06;
rommem[761] <= 16'h7C00;
rommem[762] <= 16'h3030;
rommem[763] <= 16'h7C30;
rommem[764] <= 16'h3030;
rommem[765] <= 16'h1C00;
rommem[766] <= 16'h0000;
rommem[767] <= 16'h6666;
rommem[768] <= 16'h6666;
rommem[769] <= 16'h3E00;
rommem[770] <= 16'h0000;
rommem[771] <= 16'h6666;
rommem[772] <= 16'h663C;
rommem[773] <= 16'h1800;
rommem[774] <= 16'h0000;
rommem[775] <= 16'hC6C6;
rommem[776] <= 16'hD6FE;
rommem[777] <= 16'h6C00;
rommem[778] <= 16'h0000;
rommem[779] <= 16'hC66C;
rommem[780] <= 16'h386C;
rommem[781] <= 16'hC600;
rommem[782] <= 16'h0000;
rommem[783] <= 16'h6666;
rommem[784] <= 16'h663C;
rommem[785] <= 16'h1830;
rommem[786] <= 16'h0000;
rommem[787] <= 16'h7E0C;
rommem[788] <= 16'h1830;
rommem[789] <= 16'h7E00;
rommem[790] <= 16'h0E18;
rommem[791] <= 16'h1870;
rommem[792] <= 16'h1818;
rommem[793] <= 16'h0E00;
rommem[794] <= 16'h1818;
rommem[795] <= 16'h1818;
rommem[796] <= 16'h1818;
rommem[797] <= 16'h1800;
rommem[798] <= 16'h7018;
rommem[799] <= 16'h180E;
rommem[800] <= 16'h1818;
rommem[801] <= 16'h7000;
rommem[802] <= 16'h729C;
rommem[803] <= 16'h0000;
rommem[804] <= 16'h0000;
rommem[805] <= 16'h0000;
rommem[806] <= 16'hFEFE;
rommem[807] <= 16'hFEFE;
rommem[808] <= 16'hFEFE;
rommem[809] <= 16'hFE00;
