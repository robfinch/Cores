rommem[0] <= 16'hFF40;
rommem[1] <= 16'h1000;
rommem[2] <= 16'hFFFC;
rommem[3] <= 16'h0010;
rommem[4] <= 16'h4141;
rommem[5] <= 16'h3030;
rommem[6] <= 16'h3030;
rommem[7] <= 16'h3030;
rommem[8] <= 16'h33FC;
rommem[9] <= 16'hA1A1;
rommem[10] <= 16'hFFDC;
rommem[11] <= 16'h0600;
rommem[12] <= 16'h7000;
rommem[13] <= 16'h7200;
rommem[14] <= 16'h7400;
rommem[15] <= 16'h7600;
rommem[16] <= 16'h7800;
rommem[17] <= 16'h7A00;
rommem[18] <= 16'h7C00;
rommem[19] <= 16'h7E00;
rommem[20] <= 16'h4288;
rommem[21] <= 16'h4289;
rommem[22] <= 16'h428A;
rommem[23] <= 16'h428B;
rommem[24] <= 16'h428C;
rommem[25] <= 16'h428D;
rommem[26] <= 16'h428E;
rommem[27] <= 16'h4E67;
rommem[28] <= 16'h41F9;
rommem[29] <= 16'h0000;
rommem[30] <= 16'h0000;
rommem[31] <= 16'h21C8;
rommem[32] <= 16'h0008;
rommem[33] <= 16'h41F9;
rommem[34] <= 16'hFFFC;
rommem[35] <= 16'h014C;
rommem[36] <= 16'h21C8;
rommem[37] <= 16'h0010;
rommem[38] <= 16'h41F9;
rommem[39] <= 16'hFFFC;
rommem[40] <= 16'h0132;
rommem[41] <= 16'h21C8;
rommem[42] <= 16'h0078;
rommem[43] <= 16'h41F9;
rommem[44] <= 16'h0000;
rommem[45] <= 16'h0000;
rommem[46] <= 16'h21C8;
rommem[47] <= 16'h007C;
rommem[48] <= 16'h41F9;
rommem[49] <= 16'hFFFC;
rommem[50] <= 16'h016E;
rommem[51] <= 16'h21C8;
rommem[52] <= 16'h00BC;
rommem[53] <= 16'h6100;
rommem[54] <= 16'h15BC;
rommem[55] <= 16'h33FC;
rommem[56] <= 16'hA2A2;
rommem[57] <= 16'hFFDC;
rommem[58] <= 16'h0600;
rommem[59] <= 16'h13FC;
rommem[60] <= 16'h0032;
rommem[61] <= 16'h0001;
rommem[62] <= 16'h041B;
rommem[63] <= 16'h13FC;
rommem[64] <= 16'h0025;
rommem[65] <= 16'h0001;
rommem[66] <= 16'h041A;
rommem[67] <= 16'h4239;
rommem[68] <= 16'h0001;
rommem[69] <= 16'h0419;
rommem[70] <= 16'h4239;
rommem[71] <= 16'h0001;
rommem[72] <= 16'h0418;
rommem[73] <= 16'h4279;
rommem[74] <= 16'h0001;
rommem[75] <= 16'h041C;
rommem[76] <= 16'h23FC;
rommem[77] <= 16'h0002;
rommem[78] <= 16'h0000;
rommem[79] <= 16'h0001;
rommem[80] <= 16'h0420;
rommem[81] <= 16'h4DF9;
rommem[82] <= 16'hFFDC;
rommem[83] <= 16'h0000;
rommem[84] <= 16'h426E;
rommem[85] <= 16'h0C06;
rommem[86] <= 16'h2D7C;
rommem[87] <= 16'h8888;
rommem[88] <= 16'h8888;
rommem[89] <= 16'h0C08;
rommem[90] <= 16'h2D7C;
rommem[91] <= 16'h0123;
rommem[92] <= 16'h4567;
rommem[93] <= 16'h0C0C;
rommem[94] <= 16'h6100;
rommem[95] <= 16'h0504;
rommem[96] <= 16'h6100;
rommem[97] <= 16'h0534;
rommem[98] <= 16'h6100;
rommem[99] <= 16'h056E;
rommem[100] <= 16'h6100;
rommem[101] <= 16'h03C8;
rommem[102] <= 16'h33FC;
rommem[103] <= 16'hA2A2;
rommem[104] <= 16'hFFDC;
rommem[105] <= 16'h0600;
rommem[106] <= 16'h4DF9;
rommem[107] <= 16'hFFDC;
rommem[108] <= 16'h0000;
rommem[109] <= 16'h3D7C;
rommem[110] <= 16'hFFFF;
rommem[111] <= 16'h0700;
rommem[112] <= 16'h2A7C;
rommem[113] <= 16'hFFE0;
rommem[114] <= 16'h0000;
rommem[115] <= 16'h3B7C;
rommem[116] <= 16'h4000;
rommem[117] <= 16'h0584;
rommem[118] <= 16'h6100;
rommem[119] <= 16'h13E4;
rommem[120] <= 16'h6100;
rommem[121] <= 16'h1480;
rommem[122] <= 16'h6100;
rommem[123] <= 16'h03B2;
rommem[124] <= 16'h33FC;
rommem[125] <= 16'hA3A3;
rommem[126] <= 16'hFFDC;
rommem[127] <= 16'h0600;
rommem[128] <= 16'h33FC;
rommem[129] <= 16'h7FFF;
rommem[130] <= 16'h0001;
rommem[131] <= 16'h0002;
rommem[132] <= 16'h33FC;
rommem[133] <= 16'h000F;
rommem[134] <= 16'h0001;
rommem[135] <= 16'h0004;
rommem[136] <= 16'h41F9;
rommem[137] <= 16'hFFFC;
rommem[138] <= 16'h1B9C;
rommem[139] <= 16'h7200;
rommem[140] <= 16'h7400;
rommem[141] <= 16'h6100;
rommem[142] <= 16'h05E0;
rommem[143] <= 16'h33FC;
rommem[144] <= 16'hA4A4;
rommem[145] <= 16'hFFDC;
rommem[146] <= 16'h0600;
rommem[147] <= 16'h47F9;
rommem[148] <= 16'hFFFC;
rommem[149] <= 16'h0130;
rommem[150] <= 16'h6000;
rommem[151] <= 16'h1236;
rommem[152] <= 16'h60FE;
rommem[153] <= 16'h52B9;
rommem[154] <= 16'h0001;
rommem[155] <= 16'h0430;
rommem[156] <= 16'h5279;
rommem[157] <= 16'h0001;
rommem[158] <= 16'h0434;
rommem[159] <= 16'h0279;
rommem[160] <= 16'h001F;
rommem[161] <= 16'h0001;
rommem[162] <= 16'h0434;
rommem[163] <= 16'h6702;
rommem[164] <= 16'h4E73;
rommem[165] <= 16'h4E73;
rommem[166] <= 16'h43F9;
rommem[167] <= 16'hFFFC;
rommem[168] <= 16'h015A;
rommem[169] <= 16'h4EB9;
rommem[170] <= 16'hFFFC;
rommem[171] <= 16'h03EC;
rommem[172] <= 16'h4E73;
rommem[173] <= 16'h496C;
rommem[174] <= 16'h6C65;
rommem[175] <= 16'h6761;
rommem[176] <= 16'h6C20;
rommem[177] <= 16'h696E;
rommem[178] <= 16'h7374;
rommem[179] <= 16'h7275;
rommem[180] <= 16'h6374;
rommem[181] <= 16'h696F;
rommem[182] <= 16'h6E00;
rommem[183] <= 16'h48E7;
rommem[184] <= 16'h8080;
rommem[185] <= 16'h41F9;
rommem[186] <= 16'hFFFC;
rommem[187] <= 16'h0188;
rommem[188] <= 16'hE580;
rommem[189] <= 16'h2070;
rommem[190] <= 16'h0000;
rommem[191] <= 16'h4E90;
rommem[192] <= 16'h4CDF;
rommem[193] <= 16'h0101;
rommem[194] <= 16'h4E73;
rommem[195] <= 16'hFFFF;
rommem[196] <= 16'hFFFC;
rommem[197] <= 16'h0228;
rommem[198] <= 16'hFFFC;
rommem[199] <= 16'h0228;
rommem[200] <= 16'hFFFC;
rommem[201] <= 16'h0228;
rommem[202] <= 16'hFFFC;
rommem[203] <= 16'h0228;
rommem[204] <= 16'hFFFC;
rommem[205] <= 16'h0228;
rommem[206] <= 16'hFFFC;
rommem[207] <= 16'h07FA;
rommem[208] <= 16'hFFFC;
rommem[209] <= 16'h027C;
rommem[210] <= 16'hFFFC;
rommem[211] <= 16'h07E8;
rommem[212] <= 16'hFFFC;
rommem[213] <= 16'h0228;
rommem[214] <= 16'hFFFC;
rommem[215] <= 16'h0228;
rommem[216] <= 16'hFFFC;
rommem[217] <= 16'h0228;
rommem[218] <= 16'hFFFC;
rommem[219] <= 16'h0436;
rommem[220] <= 16'hFFFC;
rommem[221] <= 16'h022A;
rommem[222] <= 16'hFFFC;
rommem[223] <= 16'h0406;
rommem[224] <= 16'hFFFC;
rommem[225] <= 16'h03EC;
rommem[226] <= 16'hFFFC;
rommem[227] <= 16'h0228;
rommem[228] <= 16'hFFFC;
rommem[229] <= 16'h0228;
rommem[230] <= 16'hFFFC;
rommem[231] <= 16'h0228;
rommem[232] <= 16'hFFFC;
rommem[233] <= 16'h0228;
rommem[234] <= 16'hFFFC;
rommem[235] <= 16'h0228;
rommem[236] <= 16'hFFFC;
rommem[237] <= 16'h0228;
rommem[238] <= 16'hFFFC;
rommem[239] <= 16'h0228;
rommem[240] <= 16'hFFFC;
rommem[241] <= 16'h0228;
rommem[242] <= 16'hFFFC;
rommem[243] <= 16'h0228;
rommem[244] <= 16'hFFFC;
rommem[245] <= 16'h0228;
rommem[246] <= 16'hFFFC;
rommem[247] <= 16'h0228;
rommem[248] <= 16'hFFFC;
rommem[249] <= 16'h0228;
rommem[250] <= 16'hFFFC;
rommem[251] <= 16'h0228;
rommem[252] <= 16'hFFFC;
rommem[253] <= 16'h0228;
rommem[254] <= 16'hFFFC;
rommem[255] <= 16'h0228;
rommem[256] <= 16'hFFFC;
rommem[257] <= 16'h0228;
rommem[258] <= 16'hFFFC;
rommem[259] <= 16'h0228;
rommem[260] <= 16'hFFFC;
rommem[261] <= 16'h0228;
rommem[262] <= 16'hFFFC;
rommem[263] <= 16'h0228;
rommem[264] <= 16'hFFFC;
rommem[265] <= 16'h0228;
rommem[266] <= 16'hFFFC;
rommem[267] <= 16'h0228;
rommem[268] <= 16'hFFFC;
rommem[269] <= 16'h0228;
rommem[270] <= 16'hFFFC;
rommem[271] <= 16'h0228;
rommem[272] <= 16'hFFFC;
rommem[273] <= 16'h0228;
rommem[274] <= 16'hFFFC;
rommem[275] <= 16'h0228;
rommem[276] <= 16'h4E75;
rommem[277] <= 16'h13C1;
rommem[278] <= 16'h0001;
rommem[279] <= 16'h0424;
rommem[280] <= 16'h4E75;
rommem[281] <= 16'h2F01;
rommem[282] <= 16'h123C;
rommem[283] <= 16'h000D;
rommem[284] <= 16'h4EB9;
rommem[285] <= 16'hFFFC;
rommem[286] <= 16'h027C;
rommem[287] <= 16'h123C;
rommem[288] <= 16'h000A;
rommem[289] <= 16'h4EB9;
rommem[290] <= 16'hFFFC;
rommem[291] <= 16'h027C;
rommem[292] <= 16'h221F;
rommem[293] <= 16'h4E75;
rommem[294] <= 16'h1039;
rommem[295] <= 16'h0001;
rommem[296] <= 16'h0418;
rommem[297] <= 16'h0240;
rommem[298] <= 16'h007F;
rommem[299] <= 16'h1439;
rommem[300] <= 16'h0001;
rommem[301] <= 16'h041B;
rommem[302] <= 16'h4882;
rommem[303] <= 16'hC0C2;
rommem[304] <= 16'h1439;
rommem[305] <= 16'h0001;
rommem[306] <= 16'h0419;
rommem[307] <= 16'h0242;
rommem[308] <= 16'h00FF;
rommem[309] <= 16'hD042;
rommem[310] <= 16'h33C0;
rommem[311] <= 16'h0001;
rommem[312] <= 16'h041C;
rommem[313] <= 16'hD0B9;
rommem[314] <= 16'h0001;
rommem[315] <= 16'h0420;
rommem[316] <= 16'h2040;
rommem[317] <= 16'h4E75;
rommem[318] <= 16'h0C01;
rommem[319] <= 16'h000D;
rommem[320] <= 16'h6608;
rommem[321] <= 16'h4239;
rommem[322] <= 16'h0001;
rommem[323] <= 16'h0419;
rommem[324] <= 16'h4E75;
rommem[325] <= 16'h0C01;
rommem[326] <= 16'h0091;
rommem[327] <= 16'h6616;
rommem[328] <= 16'h0C39;
rommem[329] <= 16'h004F;
rommem[330] <= 16'h0001;
rommem[331] <= 16'h0419;
rommem[332] <= 16'h670A;
rommem[333] <= 16'h5239;
rommem[334] <= 16'h0001;
rommem[335] <= 16'h0419;
rommem[336] <= 16'h6000;
rommem[337] <= 16'h02EA;
rommem[338] <= 16'h4E75;
rommem[339] <= 16'h0C01;
rommem[340] <= 16'h0090;
rommem[341] <= 16'h6614;
rommem[342] <= 16'h0C39;
rommem[343] <= 16'h0000;
rommem[344] <= 16'h0001;
rommem[345] <= 16'h0418;
rommem[346] <= 16'h67EE;
rommem[347] <= 16'h5339;
rommem[348] <= 16'h0001;
rommem[349] <= 16'h0418;
rommem[350] <= 16'h6000;
rommem[351] <= 16'h02CE;
rommem[352] <= 16'h0C01;
rommem[353] <= 16'h0093;
rommem[354] <= 16'h6614;
rommem[355] <= 16'h0C39;
rommem[356] <= 16'h0000;
rommem[357] <= 16'h0001;
rommem[358] <= 16'h0419;
rommem[359] <= 16'h67D4;
rommem[360] <= 16'h5339;
rommem[361] <= 16'h0001;
rommem[362] <= 16'h0419;
rommem[363] <= 16'h6000;
rommem[364] <= 16'h02B4;
rommem[365] <= 16'h0C01;
rommem[366] <= 16'h0092;
rommem[367] <= 16'h6614;
rommem[368] <= 16'h0C39;
rommem[369] <= 16'h003F;
rommem[370] <= 16'h0001;
rommem[371] <= 16'h0418;
rommem[372] <= 16'h67BA;
rommem[373] <= 16'h5279;
rommem[374] <= 16'h0001;
rommem[375] <= 16'h0418;
rommem[376] <= 16'h6000;
rommem[377] <= 16'h029A;
rommem[378] <= 16'h0C01;
rommem[379] <= 16'h0094;
rommem[380] <= 16'h661E;
rommem[381] <= 16'h0C39;
rommem[382] <= 16'h0000;
rommem[383] <= 16'h0001;
rommem[384] <= 16'h0419;
rommem[385] <= 16'h670A;
rommem[386] <= 16'h4239;
rommem[387] <= 16'h0001;
rommem[388] <= 16'h0419;
rommem[389] <= 16'h6000;
rommem[390] <= 16'h0280;
rommem[391] <= 16'h4239;
rommem[392] <= 16'h0001;
rommem[393] <= 16'h0418;
rommem[394] <= 16'h6000;
rommem[395] <= 16'h0276;
rommem[396] <= 16'h48E7;
rommem[397] <= 16'hE080;
rommem[398] <= 16'h0C01;
rommem[399] <= 16'h0099;
rommem[400] <= 16'h660C;
rommem[401] <= 16'h6100;
rommem[402] <= 16'hFF28;
rommem[403] <= 16'h1039;
rommem[404] <= 16'h0001;
rommem[405] <= 16'h0419;
rommem[406] <= 16'h6020;
rommem[407] <= 16'h0C01;
rommem[408] <= 16'h0008;
rommem[409] <= 16'h6632;
rommem[410] <= 16'h0C39;
rommem[411] <= 16'h0000;
rommem[412] <= 16'h0001;
rommem[413] <= 16'h0419;
rommem[414] <= 16'h6752;
rommem[415] <= 16'h5339;
rommem[416] <= 16'h0001;
rommem[417] <= 16'h0419;
rommem[418] <= 16'h6100;
rommem[419] <= 16'hFF06;
rommem[420] <= 16'h1039;
rommem[421] <= 16'h0001;
rommem[422] <= 16'h0419;
rommem[423] <= 16'h10E8;
rommem[424] <= 16'h0001;
rommem[425] <= 16'h5200;
rommem[426] <= 16'hB039;
rommem[427] <= 16'h0001;
rommem[428] <= 16'h041B;
rommem[429] <= 16'h65F2;
rommem[430] <= 16'h103C;
rommem[431] <= 16'h0020;
rommem[432] <= 16'h1140;
rommem[433] <= 16'hFFFF;
rommem[434] <= 16'h602A;
rommem[435] <= 16'h0C01;
rommem[436] <= 16'h000A;
rommem[437] <= 16'h671C;
rommem[438] <= 16'h6100;
rommem[439] <= 16'hFEDE;
rommem[440] <= 16'h1081;
rommem[441] <= 16'h1001;
rommem[442] <= 16'h4880;
rommem[443] <= 16'h6100;
rommem[444] <= 16'h01BA;
rommem[445] <= 16'h6100;
rommem[446] <= 16'h001A;
rommem[447] <= 16'h6100;
rommem[448] <= 16'h020C;
rommem[449] <= 16'h4CDF;
rommem[450] <= 16'h0107;
rommem[451] <= 16'h4E75;
rommem[452] <= 16'h6100;
rommem[453] <= 16'h002C;
rommem[454] <= 16'h6100;
rommem[455] <= 16'h01FE;
rommem[456] <= 16'h4CDF;
rommem[457] <= 16'h0107;
rommem[458] <= 16'h4E75;
rommem[459] <= 16'h5279;
rommem[460] <= 16'h0001;
rommem[461] <= 16'h041C;
rommem[462] <= 16'h5239;
rommem[463] <= 16'h0001;
rommem[464] <= 16'h0419;
rommem[465] <= 16'h1039;
rommem[466] <= 16'h0001;
rommem[467] <= 16'h041B;
rommem[468] <= 16'hB039;
rommem[469] <= 16'h0001;
rommem[470] <= 16'h0419;
rommem[471] <= 16'h643A;
rommem[472] <= 16'h4239;
rommem[473] <= 16'h0001;
rommem[474] <= 16'h0419;
rommem[475] <= 16'h5239;
rommem[476] <= 16'h0001;
rommem[477] <= 16'h0418;
rommem[478] <= 16'h1039;
rommem[479] <= 16'h0001;
rommem[480] <= 16'h041A;
rommem[481] <= 16'hB039;
rommem[482] <= 16'h0001;
rommem[483] <= 16'h0418;
rommem[484] <= 16'h6220;
rommem[485] <= 16'h1039;
rommem[486] <= 16'h0001;
rommem[487] <= 16'h041A;
rommem[488] <= 16'h13C0;
rommem[489] <= 16'h0001;
rommem[490] <= 16'h0418;
rommem[491] <= 16'h5339;
rommem[492] <= 16'h0001;
rommem[493] <= 16'h0418;
rommem[494] <= 16'h4880;
rommem[495] <= 16'hE340;
rommem[496] <= 16'h9179;
rommem[497] <= 16'h0001;
rommem[498] <= 16'h041C;
rommem[499] <= 16'h6100;
rommem[500] <= 16'h0CA8;
rommem[501] <= 16'h4E75;
rommem[502] <= 16'h48E7;
rommem[503] <= 16'hC040;
rommem[504] <= 16'h4281;
rommem[505] <= 16'h1219;
rommem[506] <= 16'h0C01;
rommem[507] <= 16'h0000;
rommem[508] <= 16'h6706;
rommem[509] <= 16'h6100;
rommem[510] <= 16'hFE80;
rommem[511] <= 16'h60F0;
rommem[512] <= 16'h4CDF;
rommem[513] <= 16'h0203;
rommem[514] <= 16'h4E75;
rommem[515] <= 16'h6100;
rommem[516] <= 16'hFFE4;
rommem[517] <= 16'h6000;
rommem[518] <= 16'hFE26;
rommem[519] <= 16'h48E7;
rommem[520] <= 16'hC040;
rommem[521] <= 16'h0241;
rommem[522] <= 16'h00FF;
rommem[523] <= 16'h2001;
rommem[524] <= 16'h1219;
rommem[525] <= 16'h0C01;
rommem[526] <= 16'h0000;
rommem[527] <= 16'h6708;
rommem[528] <= 16'h6100;
rommem[529] <= 16'hFE5A;
rommem[530] <= 16'h57C8;
rommem[531] <= 16'hFFF2;
rommem[532] <= 16'h4CDF;
rommem[533] <= 16'h0203;
rommem[534] <= 16'h4E75;
rommem[535] <= 16'h6100;
rommem[536] <= 16'hFFDE;
rommem[537] <= 16'h6000;
rommem[538] <= 16'hFDFE;
rommem[539] <= 16'h0C41;
rommem[540] <= 16'h00FF;
rommem[541] <= 16'h670E;
rommem[542] <= 16'h0C41;
rommem[543] <= 16'hFF00;
rommem[544] <= 16'h6718;
rommem[545] <= 16'h4EB9;
rommem[546] <= 16'hFFFC;
rommem[547] <= 16'h103E;
rommem[548] <= 16'h4E75;
rommem[549] <= 16'h1239;
rommem[550] <= 16'h0001;
rommem[551] <= 16'h0419;
rommem[552] <= 16'hE141;
rommem[553] <= 16'h1239;
rommem[554] <= 16'h0001;
rommem[555] <= 16'h0418;
rommem[556] <= 16'h4E75;
rommem[557] <= 16'h48E7;
rommem[558] <= 16'h6000;
rommem[559] <= 16'h13C1;
rommem[560] <= 16'h0001;
rommem[561] <= 16'h0418;
rommem[562] <= 16'hE049;
rommem[563] <= 16'h13C1;
rommem[564] <= 16'h0001;
rommem[565] <= 16'h0419;
rommem[566] <= 16'h1239;
rommem[567] <= 16'h0001;
rommem[568] <= 16'h0418;
rommem[569] <= 16'h4881;
rommem[570] <= 16'h1439;
rommem[571] <= 16'h0001;
rommem[572] <= 16'h041B;
rommem[573] <= 16'h4882;
rommem[574] <= 16'hC2C2;
rommem[575] <= 16'h1439;
rommem[576] <= 16'h0001;
rommem[577] <= 16'h0419;
rommem[578] <= 16'hD242;
rommem[579] <= 16'h33C1;
rommem[580] <= 16'h0001;
rommem[581] <= 16'h041C;
rommem[582] <= 16'h4CDF;
rommem[583] <= 16'h0006;
rommem[584] <= 16'h4E75;
rommem[585] <= 16'h207C;
rommem[586] <= 16'hFF80;
rommem[587] <= 16'h0000;
rommem[588] <= 16'h700F;
rommem[589] <= 16'h223C;
rommem[590] <= 16'h0001;
rommem[591] <= 16'hD4C0;
rommem[592] <= 16'h30C0;
rommem[593] <= 16'h5381;
rommem[594] <= 16'h66FA;
rommem[595] <= 16'h4E75;
rommem[596] <= 16'h2C7C;
rommem[597] <= 16'hFFE0;
rommem[598] <= 16'h0000;
rommem[599] <= 16'h2D7C;
rommem[600] <= 16'h0005;
rommem[601] <= 16'hC000;
rommem[602] <= 16'h0590;
rommem[603] <= 16'h203C;
rommem[604] <= 16'h0005;
rommem[605] <= 16'hC004;
rommem[606] <= 16'h4840;
rommem[607] <= 16'h0040;
rommem[608] <= 16'h9CE0;
rommem[609] <= 16'h4840;
rommem[610] <= 16'h23C0;
rommem[611] <= 16'hFF8B;
rommem[612] <= 16'h8000;
rommem[613] <= 16'h42B9;
rommem[614] <= 16'hFF8B;
rommem[615] <= 16'h8004;
rommem[616] <= 16'h227C;
rommem[617] <= 16'hFF8B;
rommem[618] <= 16'h8008;
rommem[619] <= 16'h41F9;
rommem[620] <= 16'hFFFC;
rommem[621] <= 16'h1C54;
rommem[622] <= 16'h223C;
rommem[623] <= 16'h0000;
rommem[624] <= 16'h1000;
rommem[625] <= 16'h3D7C;
rommem[626] <= 16'h0000;
rommem[627] <= 16'h0594;
rommem[628] <= 16'h7000;
rommem[629] <= 16'h1018;
rommem[630] <= 16'h32C0;
rommem[631] <= 16'h51C9;
rommem[632] <= 16'hFFFA;
rommem[633] <= 16'h4E75;
rommem[634] <= 16'h2C7C;
rommem[635] <= 16'hFFE0;
rommem[636] <= 16'h0000;
rommem[637] <= 16'h4840;
rommem[638] <= 16'h302E;
rommem[639] <= 16'h042C;
rommem[640] <= 16'hB07C;
rommem[641] <= 16'h001C;
rommem[642] <= 16'h64F6;
rommem[643] <= 16'h4840;
rommem[644] <= 16'h3D40;
rommem[645] <= 16'h0420;
rommem[646] <= 16'h3D79;
rommem[647] <= 16'h0001;
rommem[648] <= 16'h0002;
rommem[649] <= 16'h0422;
rommem[650] <= 16'h3D79;
rommem[651] <= 16'h0001;
rommem[652] <= 16'h0004;
rommem[653] <= 16'h0424;
rommem[654] <= 16'h3D41;
rommem[655] <= 16'h0426;
rommem[656] <= 16'h3D42;
rommem[657] <= 16'h0428;
rommem[658] <= 16'h3D7C;
rommem[659] <= 16'h0707;
rommem[660] <= 16'h042A;
rommem[661] <= 16'h3D7C;
rommem[662] <= 16'h0000;
rommem[663] <= 16'h042E;
rommem[664] <= 16'h4E75;
rommem[665] <= 16'h48E7;
rommem[666] <= 16'h4002;
rommem[667] <= 16'h2C7C;
rommem[668] <= 16'hFFE0;
rommem[669] <= 16'h0000;
rommem[670] <= 16'h4840;
rommem[671] <= 16'h302E;
rommem[672] <= 16'h042C;
rommem[673] <= 16'hB07C;
rommem[674] <= 16'h001C;
rommem[675] <= 16'h64F6;
rommem[676] <= 16'h4840;
rommem[677] <= 16'h3D40;
rommem[678] <= 16'h0420;
rommem[679] <= 16'h3D79;
rommem[680] <= 16'h0001;
rommem[681] <= 16'h0002;
rommem[682] <= 16'h0422;
rommem[683] <= 16'h3D79;
rommem[684] <= 16'h0001;
rommem[685] <= 16'h0004;
rommem[686] <= 16'h0424;
rommem[687] <= 16'h1239;
rommem[688] <= 16'h0001;
rommem[689] <= 16'h0419;
rommem[690] <= 16'h4881;
rommem[691] <= 16'hE741;
rommem[692] <= 16'h3D41;
rommem[693] <= 16'h0426;
rommem[694] <= 16'h1239;
rommem[695] <= 16'h0001;
rommem[696] <= 16'h0418;
rommem[697] <= 16'h4881;
rommem[698] <= 16'hE741;
rommem[699] <= 16'h3D41;
rommem[700] <= 16'h0428;
rommem[701] <= 16'h3D7C;
rommem[702] <= 16'h0707;
rommem[703] <= 16'h042A;
rommem[704] <= 16'h3D7C;
rommem[705] <= 16'h0000;
rommem[706] <= 16'h042E;
rommem[707] <= 16'h4CDF;
rommem[708] <= 16'h4002;
rommem[709] <= 16'h4E75;
rommem[710] <= 16'h48E7;
rommem[711] <= 16'h4002;
rommem[712] <= 16'h2C7C;
rommem[713] <= 16'hFFE0;
rommem[714] <= 16'h0000;
rommem[715] <= 16'h3D7C;
rommem[716] <= 16'h0A0A;
rommem[717] <= 16'h0444;
rommem[718] <= 16'h1239;
rommem[719] <= 16'h0001;
rommem[720] <= 16'h0419;
rommem[721] <= 16'h4881;
rommem[722] <= 16'hE741;
rommem[723] <= 16'h5341;
rommem[724] <= 16'h3D41;
rommem[725] <= 16'h0440;
rommem[726] <= 16'h1239;
rommem[727] <= 16'h0001;
rommem[728] <= 16'h0418;
rommem[729] <= 16'h4881;
rommem[730] <= 16'hE741;
rommem[731] <= 16'h5341;
rommem[732] <= 16'h3D41;
rommem[733] <= 16'h0442;
rommem[734] <= 16'h4CDF;
rommem[735] <= 16'h4002;
rommem[736] <= 16'h4E75;
rommem[737] <= 16'h2F02;
rommem[738] <= 16'h2A7C;
rommem[739] <= 16'hFFDC;
rommem[740] <= 16'h0000;
rommem[741] <= 16'h2C7C;
rommem[742] <= 16'hFFE0;
rommem[743] <= 16'h0000;
rommem[744] <= 16'h3D7C;
rommem[745] <= 16'h0004;
rommem[746] <= 16'h0446;
rommem[747] <= 16'h3D7C;
rommem[748] <= 16'h7FFF;
rommem[749] <= 16'h0448;
rommem[750] <= 16'h743F;
rommem[751] <= 16'h426D;
rommem[752] <= 16'h0C04;
rommem[753] <= 16'h262D;
rommem[754] <= 16'h0C00;
rommem[755] <= 16'h0283;
rommem[756] <= 16'h0000;
rommem[757] <= 16'hFFFF;
rommem[758] <= 16'h2CC3;
rommem[759] <= 16'h51CA;
rommem[760] <= 16'hFFEE;
rommem[761] <= 16'h241F;
rommem[762] <= 16'h4E75;
rommem[763] <= 16'h48E7;
rommem[764] <= 16'h4082;
rommem[765] <= 16'h41F9;
rommem[766] <= 16'hFFFC;
rommem[767] <= 16'h0614;
rommem[768] <= 16'h2C7C;
rommem[769] <= 16'hFFE0;
rommem[770] <= 16'h0460;
rommem[771] <= 16'h720F;
rommem[772] <= 16'h3CD8;
rommem[773] <= 16'h51C9;
rommem[774] <= 16'hFFFC;
rommem[775] <= 16'h4CDF;
rommem[776] <= 16'h4102;
rommem[777] <= 16'h4E75;
rommem[778] <= 16'h03FF;
rommem[779] <= 16'h0201;
rommem[780] <= 16'h0201;
rommem[781] <= 16'h0201;
rommem[782] <= 16'h0201;
rommem[783] <= 16'h0201;
rommem[784] <= 16'h0201;
rommem[785] <= 16'h0201;
rommem[786] <= 16'h0231;
rommem[787] <= 16'h03FF;
rommem[788] <= 16'h0000;
rommem[789] <= 16'h0000;
rommem[790] <= 16'h0000;
rommem[791] <= 16'h0000;
rommem[792] <= 16'h0000;
rommem[793] <= 16'h0000;
rommem[794] <= 16'h48E7;
rommem[795] <= 16'h70C2;
rommem[796] <= 16'h41F9;
rommem[797] <= 16'hFFFC;
rommem[798] <= 16'h069C;
rommem[799] <= 16'h7214;
rommem[800] <= 16'h227C;
rommem[801] <= 16'hFF8B;
rommem[802] <= 16'h7E00;
rommem[803] <= 16'h22D8;
rommem[804] <= 16'h51C9;
rommem[805] <= 16'hFFFC;
rommem[806] <= 16'h343C;
rommem[807] <= 16'h0200;
rommem[808] <= 16'h207C;
rommem[809] <= 16'hFFE0;
rommem[810] <= 16'h0000;
rommem[811] <= 16'h2C7C;
rommem[812] <= 16'hFFDC;
rommem[813] <= 16'h0000;
rommem[814] <= 16'h21BC;
rommem[815] <= 16'h0005;
rommem[816] <= 16'hBF00;
rommem[817] <= 16'h2000;
rommem[818] <= 16'h31BC;
rommem[819] <= 16'h0249;
rommem[820] <= 16'h2008;
rommem[821] <= 16'h426E;
rommem[822] <= 16'h0C04;
rommem[823] <= 16'h262E;
rommem[824] <= 16'h0C00;
rommem[825] <= 16'h0243;
rommem[826] <= 16'h00FF;
rommem[827] <= 16'h3183;
rommem[828] <= 16'h2004;
rommem[829] <= 16'h426E;
rommem[830] <= 16'h0C04;
rommem[831] <= 16'h262E;
rommem[832] <= 16'h0C00;
rommem[833] <= 16'h0243;
rommem[834] <= 16'h00FF;
rommem[835] <= 16'h3183;
rommem[836] <= 16'h2006;
rommem[837] <= 16'h0642;
rommem[838] <= 16'h0010;
rommem[839] <= 16'hB47C;
rommem[840] <= 16'h0300;
rommem[841] <= 16'h66C8;
rommem[842] <= 16'h4CDF;
rommem[843] <= 16'h430E;
rommem[844] <= 16'h4E75;
rommem[845] <= 16'hFFFF;
rommem[846] <= 16'h5555;
rommem[847] <= 16'h5000;
rommem[848] <= 16'h0000;
rommem[849] <= 16'h0000;
rommem[850] <= 16'h4020;
rommem[851] <= 16'h1000;
rommem[852] <= 16'h0000;
rommem[853] <= 16'h0000;
rommem[854] <= 16'h4020;
rommem[855] <= 16'h1000;
rommem[856] <= 16'h0000;
rommem[857] <= 16'h0000;
rommem[858] <= 16'h4020;
rommem[859] <= 16'h1000;
rommem[860] <= 16'h0000;
rommem[861] <= 16'h0000;
rommem[862] <= 16'h6AAA;
rommem[863] <= 16'h9000;
rommem[864] <= 16'h0000;
rommem[865] <= 16'h0000;
rommem[866] <= 16'h4020;
rommem[867] <= 16'h1000;
rommem[868] <= 16'h0000;
rommem[869] <= 16'h0000;
rommem[870] <= 16'h4020;
rommem[871] <= 16'h1000;
rommem[872] <= 16'h0000;
rommem[873] <= 16'h0000;
rommem[874] <= 16'h4020;
rommem[875] <= 16'h1000;
rommem[876] <= 16'h0000;
rommem[877] <= 16'h0000;
rommem[878] <= 16'h4050;
rommem[879] <= 16'h1000;
rommem[880] <= 16'h0000;
rommem[881] <= 16'h0000;
rommem[882] <= 16'h5555;
rommem[883] <= 16'h5000;
rommem[884] <= 16'h0000;
rommem[885] <= 16'h0000;
rommem[886] <= 16'h0000;
rommem[887] <= 16'h0000;
rommem[888] <= 16'h0000;
rommem[889] <= 16'h0000;
rommem[890] <= 16'h0000;
rommem[891] <= 16'h0000;
rommem[892] <= 16'h0000;
rommem[893] <= 16'h0000;
rommem[894] <= 16'h7000;
rommem[895] <= 16'h1018;
rommem[896] <= 16'h6708;
rommem[897] <= 16'h6100;
rommem[898] <= 16'hFDF0;
rommem[899] <= 16'h5041;
rommem[900] <= 16'h60F2;
rommem[901] <= 16'h4E75;
rommem[902] <= 16'h3F01;
rommem[903] <= 16'h0201;
rommem[904] <= 16'h000F;
rommem[905] <= 16'h0601;
rommem[906] <= 16'h0030;
rommem[907] <= 16'h0C01;
rommem[908] <= 16'h0039;
rommem[909] <= 16'h6302;
rommem[910] <= 16'h5E01;
rommem[911] <= 16'h6100;
rommem[912] <= 16'hFB5C;
rommem[913] <= 16'h321F;
rommem[914] <= 16'h4E75;
rommem[915] <= 16'h3F01;
rommem[916] <= 16'hE819;
rommem[917] <= 16'h6100;
rommem[918] <= 16'hFFE0;
rommem[919] <= 16'hE919;
rommem[920] <= 16'h6100;
rommem[921] <= 16'hFFDA;
rommem[922] <= 16'h321F;
rommem[923] <= 16'h4E75;
rommem[924] <= 16'hE199;
rommem[925] <= 16'h6100;
rommem[926] <= 16'hFFEA;
rommem[927] <= 16'hE199;
rommem[928] <= 16'h6100;
rommem[929] <= 16'hFFE4;
rommem[930] <= 16'hE199;
rommem[931] <= 16'h6100;
rommem[932] <= 16'hFFDE;
rommem[933] <= 16'hE199;
rommem[934] <= 16'h6100;
rommem[935] <= 16'hFFD8;
rommem[936] <= 16'h4E75;
rommem[937] <= 16'h123C;
rommem[938] <= 16'h003A;
rommem[939] <= 16'h4EB9;
rommem[940] <= 16'hFFFC;
rommem[941] <= 16'h027C;
rommem[942] <= 16'h2208;
rommem[943] <= 16'h4EB9;
rommem[944] <= 16'hFFFC;
rommem[945] <= 16'h0738;
rommem[946] <= 16'h7407;
rommem[947] <= 16'h123C;
rommem[948] <= 16'h0020;
rommem[949] <= 16'h4EB9;
rommem[950] <= 16'hFFFC;
rommem[951] <= 16'h027C;
rommem[952] <= 16'h1218;
rommem[953] <= 16'h4EB9;
rommem[954] <= 16'hFFFC;
rommem[955] <= 16'h0726;
rommem[956] <= 16'h51CA;
rommem[957] <= 16'hFFEC;
rommem[958] <= 16'h4EF9;
rommem[959] <= 16'hFFFC;
rommem[960] <= 16'h0232;
rommem[961] <= 16'h1239;
rommem[962] <= 16'hFFDC;
rommem[963] <= 16'h0001;
rommem[964] <= 16'h4E75;
rommem[965] <= 16'h7200;
rommem[966] <= 16'h1239;
rommem[967] <= 16'hFFDC;
rommem[968] <= 16'h0000;
rommem[969] <= 16'h13FC;
rommem[970] <= 16'h0000;
rommem[971] <= 16'hFFDC;
rommem[972] <= 16'h0001;
rommem[973] <= 16'h4E75;
rommem[974] <= 16'h2F03;
rommem[975] <= 16'h363C;
rommem[976] <= 16'h0064;
rommem[977] <= 16'h6100;
rommem[978] <= 16'hFFDE;
rommem[979] <= 16'h4A01;
rommem[980] <= 16'h6B0E;
rommem[981] <= 16'h6100;
rommem[982] <= 16'h02C4;
rommem[983] <= 16'h51CB;
rommem[984] <= 16'hFFF2;
rommem[985] <= 16'h261F;
rommem[986] <= 16'h72FF;
rommem[987] <= 16'h4E75;
rommem[988] <= 16'h6100;
rommem[989] <= 16'hFFD0;
rommem[990] <= 16'h261F;
rommem[991] <= 16'h4E75;
rommem[992] <= 16'h48E7;
rommem[993] <= 16'h3000;
rommem[994] <= 16'h7664;
rommem[995] <= 16'h6100;
rommem[996] <= 16'hFFBA;
rommem[997] <= 16'h0801;
rommem[998] <= 16'h0006;
rommem[999] <= 16'h6610;
rommem[1000] <= 16'h6100;
rommem[1001] <= 16'h029E;
rommem[1002] <= 16'h51CB;
rommem[1003] <= 16'hFFF0;
rommem[1004] <= 16'h4CDF;
rommem[1005] <= 16'h000C;
rommem[1006] <= 16'h72FF;
rommem[1007] <= 16'h4E75;
rommem[1008] <= 16'h4CDF;
rommem[1009] <= 16'h000C;
rommem[1010] <= 16'h7200;
rommem[1011] <= 16'h4E75;
rommem[1012] <= 16'h1239;
rommem[1013] <= 16'hFFDC;
rommem[1014] <= 16'h0001;
rommem[1015] <= 16'h6A06;
rommem[1016] <= 16'h123C;
rommem[1017] <= 16'h0001;
rommem[1018] <= 16'h4E75;
rommem[1019] <= 16'h4201;
rommem[1020] <= 16'h4E75;
rommem[1021] <= 16'h6100;
rommem[1022] <= 16'h0022;
rommem[1023] <= 16'h0C39;
rommem[1024] <= 16'h0000;
rommem[1025] <= 16'h0001;
rommem[1026] <= 16'h0424;
rommem[1027] <= 16'h670C;
rommem[1028] <= 16'h0C01;
rommem[1029] <= 16'h000D;
rommem[1030] <= 16'h6700;
rommem[1031] <= 16'hFA24;
rommem[1032] <= 16'h6100;
rommem[1033] <= 16'hFA6A;
rommem[1034] <= 16'h4E75;
rommem[1035] <= 16'h4239;
rommem[1036] <= 16'h0001;
rommem[1037] <= 16'h0425;
rommem[1038] <= 16'h6008;
rommem[1039] <= 16'h13FC;
rommem[1040] <= 16'hFFFF;
rommem[1041] <= 16'h0001;
rommem[1042] <= 16'h0425;
rommem[1043] <= 16'h48E7;
rommem[1044] <= 16'h3080;
rommem[1045] <= 16'h6100;
rommem[1046] <= 16'hFF56;
rommem[1047] <= 16'h6B10;
rommem[1048] <= 16'h4A39;
rommem[1049] <= 16'h0001;
rommem[1050] <= 16'h0425;
rommem[1051] <= 16'h6BF2;
rommem[1052] <= 16'h4CDF;
rommem[1053] <= 16'h010C;
rommem[1054] <= 16'h72FF;
rommem[1055] <= 16'h4E75;
rommem[1056] <= 16'h6100;
rommem[1057] <= 16'hFF48;
rommem[1058] <= 16'h33FC;
rommem[1059] <= 16'h0001;
rommem[1060] <= 16'hFFDC;
rommem[1061] <= 16'h0600;
rommem[1062] <= 16'hB23C;
rommem[1063] <= 16'h00F0;
rommem[1064] <= 16'h6700;
rommem[1065] <= 16'h00CA;
rommem[1066] <= 16'hB23C;
rommem[1067] <= 16'h00E0;
rommem[1068] <= 16'h6700;
rommem[1069] <= 16'h00CE;
rommem[1070] <= 16'hB23C;
rommem[1071] <= 16'h0014;
rommem[1072] <= 16'h6700;
rommem[1073] <= 16'h00D2;
rommem[1074] <= 16'hB23C;
rommem[1075] <= 16'h0012;
rommem[1076] <= 16'h6700;
rommem[1077] <= 16'h0134;
rommem[1078] <= 16'hB23C;
rommem[1079] <= 16'h0059;
rommem[1080] <= 16'h6700;
rommem[1081] <= 16'h012C;
rommem[1082] <= 16'hB23C;
rommem[1083] <= 16'h0077;
rommem[1084] <= 16'h6700;
rommem[1085] <= 16'h014C;
rommem[1086] <= 16'hB23C;
rommem[1087] <= 16'h0058;
rommem[1088] <= 16'h6700;
rommem[1089] <= 16'h0154;
rommem[1090] <= 16'hB23C;
rommem[1091] <= 16'h007E;
rommem[1092] <= 16'h6700;
rommem[1093] <= 16'h015C;
rommem[1094] <= 16'hB23C;
rommem[1095] <= 16'h0011;
rommem[1096] <= 16'h6700;
rommem[1097] <= 16'h00CA;
rommem[1098] <= 16'h1439;
rommem[1099] <= 16'h0001;
rommem[1100] <= 16'h0426;
rommem[1101] <= 16'h13FC;
rommem[1102] <= 16'h0000;
rommem[1103] <= 16'h0001;
rommem[1104] <= 16'h0426;
rommem[1105] <= 16'h4A02;
rommem[1106] <= 16'h6684;
rommem[1107] <= 16'hB23C;
rommem[1108] <= 16'h000D;
rommem[1109] <= 16'h6700;
rommem[1110] <= 16'h00D8;
rommem[1111] <= 16'h1439;
rommem[1112] <= 16'h0001;
rommem[1113] <= 16'h0427;
rommem[1114] <= 16'h6A1E;
rommem[1115] <= 16'h0202;
rommem[1116] <= 16'h007F;
rommem[1117] <= 16'h13C2;
rommem[1118] <= 16'h0001;
rommem[1119] <= 16'h0427;
rommem[1120] <= 16'h13FC;
rommem[1121] <= 16'h0000;
rommem[1122] <= 16'h0001;
rommem[1123] <= 16'h0426;
rommem[1124] <= 16'h41F9;
rommem[1125] <= 16'hFFFC;
rommem[1126] <= 16'h0D00;
rommem[1127] <= 16'h1230;
rommem[1128] <= 16'h1000;
rommem[1129] <= 16'h603A;
rommem[1130] <= 16'h0802;
rommem[1131] <= 16'h0002;
rommem[1132] <= 16'h6710;
rommem[1133] <= 16'h0241;
rommem[1134] <= 16'h007F;
rommem[1135] <= 16'h41F9;
rommem[1136] <= 16'hFFFC;
rommem[1137] <= 16'h0C80;
rommem[1138] <= 16'h1230;
rommem[1139] <= 16'h1000;
rommem[1140] <= 16'h6024;
rommem[1141] <= 16'h0802;
rommem[1142] <= 16'h0000;
rommem[1143] <= 16'h670C;
rommem[1144] <= 16'h41F9;
rommem[1145] <= 16'hFFFC;
rommem[1146] <= 16'h0B80;
rommem[1147] <= 16'h1230;
rommem[1148] <= 16'h1000;
rommem[1149] <= 16'h6012;
rommem[1150] <= 16'h41F9;
rommem[1151] <= 16'hFFFC;
rommem[1152] <= 16'h0A80;
rommem[1153] <= 16'h1230;
rommem[1154] <= 16'h1000;
rommem[1155] <= 16'h33FC;
rommem[1156] <= 16'h0202;
rommem[1157] <= 16'hFFDC;
rommem[1158] <= 16'h0600;
rommem[1159] <= 16'h33FC;
rommem[1160] <= 16'h0303;
rommem[1161] <= 16'hFFDC;
rommem[1162] <= 16'h0600;
rommem[1163] <= 16'h4CDF;
rommem[1164] <= 16'h010C;
rommem[1165] <= 16'h4E75;
rommem[1166] <= 16'h13FC;
rommem[1167] <= 16'hFFFF;
rommem[1168] <= 16'h0001;
rommem[1169] <= 16'h0426;
rommem[1170] <= 16'h6000;
rommem[1171] <= 16'hFF04;
rommem[1172] <= 16'h0039;
rommem[1173] <= 16'h0080;
rommem[1174] <= 16'h0001;
rommem[1175] <= 16'h0427;
rommem[1176] <= 16'h6000;
rommem[1177] <= 16'hFEF8;
rommem[1178] <= 16'h1239;
rommem[1179] <= 16'h0001;
rommem[1180] <= 16'h0426;
rommem[1181] <= 16'h4239;
rommem[1182] <= 16'h0001;
rommem[1183] <= 16'h0426;
rommem[1184] <= 16'h4A01;
rommem[1185] <= 16'h6A0C;
rommem[1186] <= 16'h08B9;
rommem[1187] <= 16'h0002;
rommem[1188] <= 16'h0001;
rommem[1189] <= 16'h0427;
rommem[1190] <= 16'h6000;
rommem[1191] <= 16'hFEDC;
rommem[1192] <= 16'h08F9;
rommem[1193] <= 16'h0002;
rommem[1194] <= 16'h0001;
rommem[1195] <= 16'h0427;
rommem[1196] <= 16'h6000;
rommem[1197] <= 16'hFED0;
rommem[1198] <= 16'h1239;
rommem[1199] <= 16'h0001;
rommem[1200] <= 16'h0426;
rommem[1201] <= 16'h4239;
rommem[1202] <= 16'h0001;
rommem[1203] <= 16'h0426;
rommem[1204] <= 16'h4A01;
rommem[1205] <= 16'h6A0C;
rommem[1206] <= 16'h08B9;
rommem[1207] <= 16'h0001;
rommem[1208] <= 16'h0001;
rommem[1209] <= 16'h0427;
rommem[1210] <= 16'h6000;
rommem[1211] <= 16'hFEB4;
rommem[1212] <= 16'h08F9;
rommem[1213] <= 16'h0001;
rommem[1214] <= 16'h0001;
rommem[1215] <= 16'h0427;
rommem[1216] <= 16'h6000;
rommem[1217] <= 16'hFEA8;
rommem[1218] <= 16'h2F01;
rommem[1219] <= 16'h1239;
rommem[1220] <= 16'h0001;
rommem[1221] <= 16'h0427;
rommem[1222] <= 16'h0801;
rommem[1223] <= 16'h0000;
rommem[1224] <= 16'h6706;
rommem[1225] <= 16'h221F;
rommem[1226] <= 16'h6000;
rommem[1227] <= 16'hFE94;
rommem[1228] <= 16'h221F;
rommem[1229] <= 16'h6000;
rommem[1230] <= 16'hFF12;
rommem[1231] <= 16'h1239;
rommem[1232] <= 16'h0001;
rommem[1233] <= 16'h0426;
rommem[1234] <= 16'h4239;
rommem[1235] <= 16'h0001;
rommem[1236] <= 16'h0426;
rommem[1237] <= 16'h4A01;
rommem[1238] <= 16'h6A0C;
rommem[1239] <= 16'h08B9;
rommem[1240] <= 16'h0000;
rommem[1241] <= 16'h0001;
rommem[1242] <= 16'h0427;
rommem[1243] <= 16'h6000;
rommem[1244] <= 16'hFE72;
rommem[1245] <= 16'h08F9;
rommem[1246] <= 16'h0000;
rommem[1247] <= 16'h0001;
rommem[1248] <= 16'h0427;
rommem[1249] <= 16'h6000;
rommem[1250] <= 16'hFE66;
rommem[1251] <= 16'h0879;
rommem[1252] <= 16'h0004;
rommem[1253] <= 16'h0001;
rommem[1254] <= 16'h0427;
rommem[1255] <= 16'h6100;
rommem[1256] <= 16'h0026;
rommem[1257] <= 16'h6000;
rommem[1258] <= 16'hFE56;
rommem[1259] <= 16'h0879;
rommem[1260] <= 16'h0005;
rommem[1261] <= 16'h0001;
rommem[1262] <= 16'h0427;
rommem[1263] <= 16'h6100;
rommem[1264] <= 16'h0016;
rommem[1265] <= 16'h6000;
rommem[1266] <= 16'hFE46;
rommem[1267] <= 16'h0879;
rommem[1268] <= 16'h0006;
rommem[1269] <= 16'h0001;
rommem[1270] <= 16'h0427;
rommem[1271] <= 16'h6100;
rommem[1272] <= 16'h0006;
rommem[1273] <= 16'h6000;
rommem[1274] <= 16'hFE36;
rommem[1275] <= 16'h48E7;
rommem[1276] <= 16'h3000;
rommem[1277] <= 16'h4239;
rommem[1278] <= 16'h0001;
rommem[1279] <= 16'h0428;
rommem[1280] <= 16'h0839;
rommem[1281] <= 16'h0004;
rommem[1282] <= 16'h0001;
rommem[1283] <= 16'h0427;
rommem[1284] <= 16'h6708;
rommem[1285] <= 16'h13FC;
rommem[1286] <= 16'h0002;
rommem[1287] <= 16'h0001;
rommem[1288] <= 16'h0428;
rommem[1289] <= 16'h0839;
rommem[1290] <= 16'h0005;
rommem[1291] <= 16'h0001;
rommem[1292] <= 16'h0427;
rommem[1293] <= 16'h6708;
rommem[1294] <= 16'h08F9;
rommem[1295] <= 16'h0002;
rommem[1296] <= 16'h0001;
rommem[1297] <= 16'h0428;
rommem[1298] <= 16'h0839;
rommem[1299] <= 16'h0006;
rommem[1300] <= 16'h0001;
rommem[1301] <= 16'h0427;
rommem[1302] <= 16'h6708;
rommem[1303] <= 16'h08F9;
rommem[1304] <= 16'h0000;
rommem[1305] <= 16'h0001;
rommem[1306] <= 16'h0428;
rommem[1307] <= 16'h123C;
rommem[1308] <= 16'h00ED;
rommem[1309] <= 16'h6100;
rommem[1310] <= 16'h002C;
rommem[1311] <= 16'h6100;
rommem[1312] <= 16'hFD80;
rommem[1313] <= 16'h6100;
rommem[1314] <= 16'hFD58;
rommem[1315] <= 16'h4A01;
rommem[1316] <= 16'h6B18;
rommem[1317] <= 16'hB2BC;
rommem[1318] <= 16'h0000;
rommem[1319] <= 16'h00FA;
rommem[1320] <= 16'h1239;
rommem[1321] <= 16'h0001;
rommem[1322] <= 16'h0428;
rommem[1323] <= 16'h6100;
rommem[1324] <= 16'h0010;
rommem[1325] <= 16'h6100;
rommem[1326] <= 16'hFD64;
rommem[1327] <= 16'h6100;
rommem[1328] <= 16'hFD3C;
rommem[1329] <= 16'h4CDF;
rommem[1330] <= 16'h000C;
rommem[1331] <= 16'h4E75;
rommem[1332] <= 16'h13C1;
rommem[1333] <= 16'hFFDC;
rommem[1334] <= 16'h0000;
rommem[1335] <= 16'h4E75;
rommem[1336] <= 16'h2F03;
rommem[1337] <= 16'h263C;
rommem[1338] <= 16'h0000;
rommem[1339] <= 16'h03E8;
rommem[1340] <= 16'h51CB;
rommem[1341] <= 16'hFFFE;
rommem[1342] <= 16'h261F;
rommem[1343] <= 16'h4E75;
rommem[1344] <= 16'h2EA9;
rommem[1345] <= 16'h2EA5;
rommem[1346] <= 16'hA3A1;
rommem[1347] <= 16'hA2AC;
rommem[1348] <= 16'h2EAA;
rommem[1349] <= 16'hA8A6;
rommem[1350] <= 16'hA409;
rommem[1351] <= 16'h602E;
rommem[1352] <= 16'h2E2E;
rommem[1353] <= 16'h2E2E;
rommem[1354] <= 16'h2E71;
rommem[1355] <= 16'h312E;
rommem[1356] <= 16'h2E2E;
rommem[1357] <= 16'h7A73;
rommem[1358] <= 16'h6177;
rommem[1359] <= 16'h322E;
rommem[1360] <= 16'h2E63;
rommem[1361] <= 16'h7864;
rommem[1362] <= 16'h6534;
rommem[1363] <= 16'h332E;
rommem[1364] <= 16'h2E20;
rommem[1365] <= 16'h7666;
rommem[1366] <= 16'h7472;
rommem[1367] <= 16'h352E;
rommem[1368] <= 16'h2E6E;
rommem[1369] <= 16'h6268;
rommem[1370] <= 16'h6779;
rommem[1371] <= 16'h362E;
rommem[1372] <= 16'h2E2E;
rommem[1373] <= 16'h6D6A;
rommem[1374] <= 16'h7537;
rommem[1375] <= 16'h382E;
rommem[1376] <= 16'h2E2C;
rommem[1377] <= 16'h6B69;
rommem[1378] <= 16'h6F30;
rommem[1379] <= 16'h392E;
rommem[1380] <= 16'h2E2E;
rommem[1381] <= 16'h2F6C;
rommem[1382] <= 16'h3B70;
rommem[1383] <= 16'h2D2E;
rommem[1384] <= 16'h2E2E;
rommem[1385] <= 16'h272E;
rommem[1386] <= 16'h5B3D;
rommem[1387] <= 16'h2E2E;
rommem[1388] <= 16'hAD2E;
rommem[1389] <= 16'h0D5D;
rommem[1390] <= 16'h2E5C;
rommem[1391] <= 16'h2E2E;
rommem[1392] <= 16'h2E2E;
rommem[1393] <= 16'h2E2E;
rommem[1394] <= 16'h2E2E;
rommem[1395] <= 16'h082E;
rommem[1396] <= 16'h2E95;
rommem[1397] <= 16'h2E93;
rommem[1398] <= 16'h942E;
rommem[1399] <= 16'h2E2E;
rommem[1400] <= 16'h987F;
rommem[1401] <= 16'h922E;
rommem[1402] <= 16'h9190;
rommem[1403] <= 16'h1BAF;
rommem[1404] <= 16'hAB2E;
rommem[1405] <= 16'h972E;
rommem[1406] <= 16'h2E96;
rommem[1407] <= 16'hAE2E;
rommem[1408] <= 16'h2E2E;
rommem[1409] <= 16'h2EA7;
rommem[1410] <= 16'h2E2E;
rommem[1411] <= 16'h2E2E;
rommem[1412] <= 16'h2E2E;
rommem[1413] <= 16'h2E2E;
rommem[1414] <= 16'h2E2E;
rommem[1415] <= 16'h2E2E;
rommem[1416] <= 16'h2E2E;
rommem[1417] <= 16'h2E2E;
rommem[1418] <= 16'h2E2E;
rommem[1419] <= 16'h2E2E;
rommem[1420] <= 16'h2E2E;
rommem[1421] <= 16'h2E2E;
rommem[1422] <= 16'h2E2E;
rommem[1423] <= 16'h2E2E;
rommem[1424] <= 16'h2E2E;
rommem[1425] <= 16'h2E2E;
rommem[1426] <= 16'h2E2E;
rommem[1427] <= 16'h2E2E;
rommem[1428] <= 16'h2E2E;
rommem[1429] <= 16'h2E2E;
rommem[1430] <= 16'h2E2E;
rommem[1431] <= 16'h2E2E;
rommem[1432] <= 16'h2E2E;
rommem[1433] <= 16'h2E2E;
rommem[1434] <= 16'h2E2E;
rommem[1435] <= 16'h2E2E;
rommem[1436] <= 16'h2E2E;
rommem[1437] <= 16'h2E2E;
rommem[1438] <= 16'h2E2E;
rommem[1439] <= 16'h2E2E;
rommem[1440] <= 16'h2E2E;
rommem[1441] <= 16'h2E2E;
rommem[1442] <= 16'h2E2E;
rommem[1443] <= 16'h2E2E;
rommem[1444] <= 16'h2E2E;
rommem[1445] <= 16'h2E2E;
rommem[1446] <= 16'h2E2E;
rommem[1447] <= 16'h2E2E;
rommem[1448] <= 16'h2E2E;
rommem[1449] <= 16'h2E2E;
rommem[1450] <= 16'h2E2E;
rommem[1451] <= 16'h2E2E;
rommem[1452] <= 16'h2E2E;
rommem[1453] <= 16'h2E2E;
rommem[1454] <= 16'h2E2E;
rommem[1455] <= 16'h2E2E;
rommem[1456] <= 16'h2E2E;
rommem[1457] <= 16'h2E2E;
rommem[1458] <= 16'h2E2E;
rommem[1459] <= 16'h2E2E;
rommem[1460] <= 16'h2E2E;
rommem[1461] <= 16'h2E2E;
rommem[1462] <= 16'h2E2E;
rommem[1463] <= 16'h2E2E;
rommem[1464] <= 16'h2E2E;
rommem[1465] <= 16'h2E2E;
rommem[1466] <= 16'h2E2E;
rommem[1467] <= 16'h2E2E;
rommem[1468] <= 16'h2E2E;
rommem[1469] <= 16'hFA2E;
rommem[1470] <= 16'h2E2E;
rommem[1471] <= 16'h2E2E;
rommem[1472] <= 16'h2E2E;
rommem[1473] <= 16'h2E2E;
rommem[1474] <= 16'h2E2E;
rommem[1475] <= 16'h2E2E;
rommem[1476] <= 16'h2E2E;
rommem[1477] <= 16'h2E2E;
rommem[1478] <= 16'h2E09;
rommem[1479] <= 16'h7E2E;
rommem[1480] <= 16'h2E2E;
rommem[1481] <= 16'h2E2E;
rommem[1482] <= 16'h2E51;
rommem[1483] <= 16'h212E;
rommem[1484] <= 16'h2E2E;
rommem[1485] <= 16'h5A53;
rommem[1486] <= 16'h4157;
rommem[1487] <= 16'h402E;
rommem[1488] <= 16'h2E43;
rommem[1489] <= 16'h5844;
rommem[1490] <= 16'h4524;
rommem[1491] <= 16'h232E;
rommem[1492] <= 16'h2E20;
rommem[1493] <= 16'h5646;
rommem[1494] <= 16'h5452;
rommem[1495] <= 16'h252E;
rommem[1496] <= 16'h2E4E;
rommem[1497] <= 16'h4248;
rommem[1498] <= 16'h4759;
rommem[1499] <= 16'h5E2E;
rommem[1500] <= 16'h2E2E;
rommem[1501] <= 16'h4D4A;
rommem[1502] <= 16'h5526;
rommem[1503] <= 16'h2A2E;
rommem[1504] <= 16'h2E3C;
rommem[1505] <= 16'h4B49;
rommem[1506] <= 16'h4F29;
rommem[1507] <= 16'h282E;
rommem[1508] <= 16'h2E3E;
rommem[1509] <= 16'h3F4C;
rommem[1510] <= 16'h3A50;
rommem[1511] <= 16'h5F2E;
rommem[1512] <= 16'h2E2E;
rommem[1513] <= 16'h222E;
rommem[1514] <= 16'h7B2B;
rommem[1515] <= 16'h2E2E;
rommem[1516] <= 16'h2E2E;
rommem[1517] <= 16'h0D7D;
rommem[1518] <= 16'h2E7C;
rommem[1519] <= 16'h2E2E;
rommem[1520] <= 16'h2E2E;
rommem[1521] <= 16'h2E2E;
rommem[1522] <= 16'h2E2E;
rommem[1523] <= 16'h082E;
rommem[1524] <= 16'h2E2E;
rommem[1525] <= 16'h2E2E;
rommem[1526] <= 16'h2E2E;
rommem[1527] <= 16'h2E2E;
rommem[1528] <= 16'h2E7F;
rommem[1529] <= 16'h2E2E;
rommem[1530] <= 16'h2E2E;
rommem[1531] <= 16'h1B2E;
rommem[1532] <= 16'h2E2E;
rommem[1533] <= 16'h2E2E;
rommem[1534] <= 16'h2E2E;
rommem[1535] <= 16'h2E2E;
rommem[1536] <= 16'h2E2E;
rommem[1537] <= 16'h2E2E;
rommem[1538] <= 16'h2E2E;
rommem[1539] <= 16'h2E2E;
rommem[1540] <= 16'h2E2E;
rommem[1541] <= 16'h2E2E;
rommem[1542] <= 16'h2E2E;
rommem[1543] <= 16'h2E2E;
rommem[1544] <= 16'h2E2E;
rommem[1545] <= 16'h2E2E;
rommem[1546] <= 16'h2E2E;
rommem[1547] <= 16'h2E2E;
rommem[1548] <= 16'h2E2E;
rommem[1549] <= 16'h2E2E;
rommem[1550] <= 16'h2E2E;
rommem[1551] <= 16'h2E2E;
rommem[1552] <= 16'h2E2E;
rommem[1553] <= 16'h2E2E;
rommem[1554] <= 16'h2E2E;
rommem[1555] <= 16'h2E2E;
rommem[1556] <= 16'h2E2E;
rommem[1557] <= 16'h2E2E;
rommem[1558] <= 16'h2E2E;
rommem[1559] <= 16'h2E2E;
rommem[1560] <= 16'h2E2E;
rommem[1561] <= 16'h2E2E;
rommem[1562] <= 16'h2E2E;
rommem[1563] <= 16'h2E2E;
rommem[1564] <= 16'h2E2E;
rommem[1565] <= 16'h2E2E;
rommem[1566] <= 16'h2E2E;
rommem[1567] <= 16'h2E2E;
rommem[1568] <= 16'h2E2E;
rommem[1569] <= 16'h2E2E;
rommem[1570] <= 16'h2E2E;
rommem[1571] <= 16'h2E2E;
rommem[1572] <= 16'h2E2E;
rommem[1573] <= 16'h2E2E;
rommem[1574] <= 16'h2E2E;
rommem[1575] <= 16'h2E2E;
rommem[1576] <= 16'h2E2E;
rommem[1577] <= 16'h2E2E;
rommem[1578] <= 16'h2E2E;
rommem[1579] <= 16'h2E2E;
rommem[1580] <= 16'h2E2E;
rommem[1581] <= 16'h2E2E;
rommem[1582] <= 16'h2E2E;
rommem[1583] <= 16'h2E2E;
rommem[1584] <= 16'h2E2E;
rommem[1585] <= 16'h2E2E;
rommem[1586] <= 16'h2E2E;
rommem[1587] <= 16'h2E2E;
rommem[1588] <= 16'h2E2E;
rommem[1589] <= 16'h2E2E;
rommem[1590] <= 16'h2E2E;
rommem[1591] <= 16'h2E2E;
rommem[1592] <= 16'h2E2E;
rommem[1593] <= 16'h2E2E;
rommem[1594] <= 16'h2E2E;
rommem[1595] <= 16'h2E2E;
rommem[1596] <= 16'h2E2E;
rommem[1597] <= 16'h2E2E;
rommem[1598] <= 16'h2E2E;
rommem[1599] <= 16'h2E2E;
rommem[1600] <= 16'h2E2E;
rommem[1601] <= 16'h2E2E;
rommem[1602] <= 16'h2E2E;
rommem[1603] <= 16'h2E2E;
rommem[1604] <= 16'h2E2E;
rommem[1605] <= 16'h2E2E;
rommem[1606] <= 16'h2E09;
rommem[1607] <= 16'h7E2E;
rommem[1608] <= 16'h2E2E;
rommem[1609] <= 16'h2E2E;
rommem[1610] <= 16'h2E11;
rommem[1611] <= 16'h212E;
rommem[1612] <= 16'h2E2E;
rommem[1613] <= 16'h1A13;
rommem[1614] <= 16'h0117;
rommem[1615] <= 16'h402E;
rommem[1616] <= 16'h2E03;
rommem[1617] <= 16'h1804;
rommem[1618] <= 16'h0524;
rommem[1619] <= 16'h232E;
rommem[1620] <= 16'h2E20;
rommem[1621] <= 16'h1606;
rommem[1622] <= 16'h1412;
rommem[1623] <= 16'h252E;
rommem[1624] <= 16'h2E0E;
rommem[1625] <= 16'h0208;
rommem[1626] <= 16'h0719;
rommem[1627] <= 16'h5E2E;
rommem[1628] <= 16'h2E2E;
rommem[1629] <= 16'h0D0A;
rommem[1630] <= 16'h1526;
rommem[1631] <= 16'h2A2E;
rommem[1632] <= 16'h2E3C;
rommem[1633] <= 16'h0B09;
rommem[1634] <= 16'h0F29;
rommem[1635] <= 16'h282E;
rommem[1636] <= 16'h2E3E;
rommem[1637] <= 16'h3F0C;
rommem[1638] <= 16'h3A10;
rommem[1639] <= 16'h5F2E;
rommem[1640] <= 16'h2E2E;
rommem[1641] <= 16'h222E;
rommem[1642] <= 16'h7B2B;
rommem[1643] <= 16'h2E2E;
rommem[1644] <= 16'h2E2E;
rommem[1645] <= 16'h0D7D;
rommem[1646] <= 16'h2E7C;
rommem[1647] <= 16'h2E2E;
rommem[1648] <= 16'h2E2E;
rommem[1649] <= 16'h2E2E;
rommem[1650] <= 16'h2E2E;
rommem[1651] <= 16'h082E;
rommem[1652] <= 16'h2E2E;
rommem[1653] <= 16'h2E2E;
rommem[1654] <= 16'h2E2E;
rommem[1655] <= 16'h2E2E;
rommem[1656] <= 16'h2E7F;
rommem[1657] <= 16'h2E2E;
rommem[1658] <= 16'h2E2E;
rommem[1659] <= 16'h1B2E;
rommem[1660] <= 16'h2E2E;
rommem[1661] <= 16'h2E2E;
rommem[1662] <= 16'h2E2E;
rommem[1663] <= 16'h2E2E;
rommem[1664] <= 16'h2E2E;
rommem[1665] <= 16'h2E2E;
rommem[1666] <= 16'hA3A1;
rommem[1667] <= 16'hA22E;
rommem[1668] <= 16'h2E2E;
rommem[1669] <= 16'h2E2E;
rommem[1670] <= 16'h2E2E;
rommem[1671] <= 16'h2E2E;
rommem[1672] <= 16'h2E2E;
rommem[1673] <= 16'h2E2E;
rommem[1674] <= 16'h2E2E;
rommem[1675] <= 16'h2E2E;
rommem[1676] <= 16'h2E2E;
rommem[1677] <= 16'h2E2E;
rommem[1678] <= 16'h2E2E;
rommem[1679] <= 16'h2E2E;
rommem[1680] <= 16'h2E2E;
rommem[1681] <= 16'h2E2E;
rommem[1682] <= 16'h2E2E;
rommem[1683] <= 16'h2E2E;
rommem[1684] <= 16'h2E2E;
rommem[1685] <= 16'h2E2E;
rommem[1686] <= 16'h2E2E;
rommem[1687] <= 16'h2E2E;
rommem[1688] <= 16'h2E2E;
rommem[1689] <= 16'h2E2E;
rommem[1690] <= 16'h2E2E;
rommem[1691] <= 16'h2E2E;
rommem[1692] <= 16'h2E2E;
rommem[1693] <= 16'h2E2E;
rommem[1694] <= 16'h2E2E;
rommem[1695] <= 16'h2E2E;
rommem[1696] <= 16'h2E2E;
rommem[1697] <= 16'h2E2E;
rommem[1698] <= 16'h2E2E;
rommem[1699] <= 16'h2E2E;
rommem[1700] <= 16'h2E2E;
rommem[1701] <= 16'h2E2E;
rommem[1702] <= 16'h2E2E;
rommem[1703] <= 16'h2E2E;
rommem[1704] <= 16'h2E2E;
rommem[1705] <= 16'h2E2E;
rommem[1706] <= 16'h2E2E;
rommem[1707] <= 16'h2E2E;
rommem[1708] <= 16'h2E2E;
rommem[1709] <= 16'h2E2E;
rommem[1710] <= 16'h2E2E;
rommem[1711] <= 16'h2E2E;
rommem[1712] <= 16'h2E2E;
rommem[1713] <= 16'h2E2E;
rommem[1714] <= 16'h2E2E;
rommem[1715] <= 16'h2E2E;
rommem[1716] <= 16'h2E95;
rommem[1717] <= 16'h2E93;
rommem[1718] <= 16'h942E;
rommem[1719] <= 16'h2E2E;
rommem[1720] <= 16'h9899;
rommem[1721] <= 16'h922E;
rommem[1722] <= 16'h9190;
rommem[1723] <= 16'h2E2E;
rommem[1724] <= 16'h2E2E;
rommem[1725] <= 16'h972E;
rommem[1726] <= 16'h2E96;
rommem[1727] <= 16'h2E2E;
rommem[1728] <= 16'h4239;
rommem[1729] <= 16'h0001;
rommem[1730] <= 16'h0424;
rommem[1731] <= 16'h6100;
rommem[1732] <= 16'hF4AA;
rommem[1733] <= 16'h123C;
rommem[1734] <= 16'h0024;
rommem[1735] <= 16'h6100;
rommem[1736] <= 16'hF4EC;
rommem[1737] <= 16'h6100;
rommem[1738] <= 16'hFA66;
rommem[1739] <= 16'h0C01;
rommem[1740] <= 16'h000D;
rommem[1741] <= 16'h6706;
rommem[1742] <= 16'h6100;
rommem[1743] <= 16'hF4DE;
rommem[1744] <= 16'h60F0;
rommem[1745] <= 16'h4239;
rommem[1746] <= 16'h0001;
rommem[1747] <= 16'h0419;
rommem[1748] <= 16'h6100;
rommem[1749] <= 16'hF4A2;
rommem[1750] <= 16'h1218;
rommem[1751] <= 16'h0C01;
rommem[1752] <= 16'h0024;
rommem[1753] <= 16'h6602;
rommem[1754] <= 16'h1218;
rommem[1755] <= 16'h0C01;
rommem[1756] <= 16'h006F;
rommem[1757] <= 16'h6700;
rommem[1758] <= 16'h0D8E;
rommem[1759] <= 16'h0C01;
rommem[1760] <= 16'h0061;
rommem[1761] <= 16'h6700;
rommem[1762] <= 16'h08DC;
rommem[1763] <= 16'h0C01;
rommem[1764] <= 16'h0067;
rommem[1765] <= 16'h6700;
rommem[1766] <= 16'h0684;
rommem[1767] <= 16'h0C01;
rommem[1768] <= 16'h003A;
rommem[1769] <= 16'h6700;
rommem[1770] <= 16'h015C;
rommem[1771] <= 16'h0C01;
rommem[1772] <= 16'h0044;
rommem[1773] <= 16'h6700;
rommem[1774] <= 16'h01C2;
rommem[1775] <= 16'h0C01;
rommem[1776] <= 16'h0046;
rommem[1777] <= 16'h6700;
rommem[1778] <= 16'h00F6;
rommem[1779] <= 16'h0C01;
rommem[1780] <= 16'h0042;
rommem[1781] <= 16'h6606;
rommem[1782] <= 16'h4EF9;
rommem[1783] <= 16'hFFFC;
rommem[1784] <= 16'hC000;
rommem[1785] <= 16'h0C01;
rommem[1786] <= 16'h004A;
rommem[1787] <= 16'h6700;
rommem[1788] <= 16'h0196;
rommem[1789] <= 16'h0C01;
rommem[1790] <= 16'h004C;
rommem[1791] <= 16'h6700;
rommem[1792] <= 16'h0368;
rommem[1793] <= 16'h0C01;
rommem[1794] <= 16'h003F;
rommem[1795] <= 16'h6726;
rommem[1796] <= 16'h0C01;
rommem[1797] <= 16'h0043;
rommem[1798] <= 16'h6704;
rommem[1799] <= 16'h6000;
rommem[1800] <= 16'hFF70;
rommem[1801] <= 16'h1218;
rommem[1802] <= 16'h0C01;
rommem[1803] <= 16'h004C;
rommem[1804] <= 16'h6600;
rommem[1805] <= 16'hFF66;
rommem[1806] <= 16'h1218;
rommem[1807] <= 16'h0C01;
rommem[1808] <= 16'h0053;
rommem[1809] <= 16'h6600;
rommem[1810] <= 16'hFF5C;
rommem[1811] <= 16'h6100;
rommem[1812] <= 16'h0216;
rommem[1813] <= 16'h6000;
rommem[1814] <= 16'hFF54;
rommem[1815] <= 16'h43F9;
rommem[1816] <= 16'hFFFC;
rommem[1817] <= 16'h0E3E;
rommem[1818] <= 16'h4EB9;
rommem[1819] <= 16'hFFFC;
rommem[1820] <= 16'h03EC;
rommem[1821] <= 16'h6000;
rommem[1822] <= 16'hFF44;
rommem[1823] <= 16'h3F20;
rommem[1824] <= 16'h3D20;
rommem[1825] <= 16'h4469;
rommem[1826] <= 16'h7370;
rommem[1827] <= 16'h6C61;
rommem[1828] <= 16'h7920;
rommem[1829] <= 16'h6865;
rommem[1830] <= 16'h6C70;
rommem[1831] <= 16'h0D0A;
rommem[1832] <= 16'h434C;
rommem[1833] <= 16'h5320;
rommem[1834] <= 16'h3D20;
rommem[1835] <= 16'h636C;
rommem[1836] <= 16'h6561;
rommem[1837] <= 16'h7220;
rommem[1838] <= 16'h7363;
rommem[1839] <= 16'h7265;
rommem[1840] <= 16'h656E;
rommem[1841] <= 16'h0D0A;
rommem[1842] <= 16'h3A20;
rommem[1843] <= 16'h3D20;
rommem[1844] <= 16'h4564;
rommem[1845] <= 16'h6974;
rommem[1846] <= 16'h206D;
rommem[1847] <= 16'h656D;
rommem[1848] <= 16'h6F72;
rommem[1849] <= 16'h7920;
rommem[1850] <= 16'h6279;
rommem[1851] <= 16'h7465;
rommem[1852] <= 16'h730D;
rommem[1853] <= 16'h0A46;
rommem[1854] <= 16'h203D;
rommem[1855] <= 16'h2046;
rommem[1856] <= 16'h696C;
rommem[1857] <= 16'h6C20;
rommem[1858] <= 16'h6D65;
rommem[1859] <= 16'h6D6F;
rommem[1860] <= 16'h7279;
rommem[1861] <= 16'h0D0A;
rommem[1862] <= 16'h4C20;
rommem[1863] <= 16'h3D20;
rommem[1864] <= 16'h4C6F;
rommem[1865] <= 16'h6164;
rommem[1866] <= 16'h2053;
rommem[1867] <= 16'h3139;
rommem[1868] <= 16'h2066;
rommem[1869] <= 16'h696C;
rommem[1870] <= 16'h650D;
rommem[1871] <= 16'h0A44;
rommem[1872] <= 16'h203D;
rommem[1873] <= 16'h2044;
rommem[1874] <= 16'h756D;
rommem[1875] <= 16'h7020;
rommem[1876] <= 16'h6D65;
rommem[1877] <= 16'h6D6F;
rommem[1878] <= 16'h7279;
rommem[1879] <= 16'h0D0A;
rommem[1880] <= 16'h4220;
rommem[1881] <= 16'h3D20;
rommem[1882] <= 16'h7374;
rommem[1883] <= 16'h6172;
rommem[1884] <= 16'h7420;
rommem[1885] <= 16'h7469;
rommem[1886] <= 16'h6E79;
rommem[1887] <= 16'h2062;
rommem[1888] <= 16'h6173;
rommem[1889] <= 16'h6963;
rommem[1890] <= 16'h0D0A;
rommem[1891] <= 16'h4A20;
rommem[1892] <= 16'h3D20;
rommem[1893] <= 16'h4A75;
rommem[1894] <= 16'h6D70;
rommem[1895] <= 16'h2074;
rommem[1896] <= 16'h6F20;
rommem[1897] <= 16'h636F;
rommem[1898] <= 16'h6465;
rommem[1899] <= 16'h0D0A;
rommem[1900] <= 16'h00FF;
rommem[1901] <= 16'h1218;
rommem[1902] <= 16'h1801;
rommem[1903] <= 16'h6100;
rommem[1904] <= 16'h0044;
rommem[1905] <= 16'h6100;
rommem[1906] <= 16'h00EE;
rommem[1907] <= 16'h2241;
rommem[1908] <= 16'h6100;
rommem[1909] <= 16'h003A;
rommem[1910] <= 16'h6100;
rommem[1911] <= 16'h00E4;
rommem[1912] <= 16'h2601;
rommem[1913] <= 16'h6100;
rommem[1914] <= 16'h0030;
rommem[1915] <= 16'h6100;
rommem[1916] <= 16'h00DA;
rommem[1917] <= 16'h0C04;
rommem[1918] <= 16'h004C;
rommem[1919] <= 16'h660A;
rommem[1920] <= 16'h22C1;
rommem[1921] <= 16'h5383;
rommem[1922] <= 16'h66FA;
rommem[1923] <= 16'h6000;
rommem[1924] <= 16'hFE78;
rommem[1925] <= 16'h0C04;
rommem[1926] <= 16'h0057;
rommem[1927] <= 16'h660A;
rommem[1928] <= 16'h32C1;
rommem[1929] <= 16'h5383;
rommem[1930] <= 16'h66FA;
rommem[1931] <= 16'h6000;
rommem[1932] <= 16'hFE68;
rommem[1933] <= 16'h12C1;
rommem[1934] <= 16'h5383;
rommem[1935] <= 16'h66FA;
rommem[1936] <= 16'h6000;
rommem[1937] <= 16'hFE5E;
rommem[1938] <= 16'h1218;
rommem[1939] <= 16'h0C01;
rommem[1940] <= 16'h0020;
rommem[1941] <= 16'h67F8;
rommem[1942] <= 16'h5388;
rommem[1943] <= 16'h4E75;
rommem[1944] <= 16'h6100;
rommem[1945] <= 16'hFFF2;
rommem[1946] <= 16'h6100;
rommem[1947] <= 16'h009C;
rommem[1948] <= 16'h2241;
rommem[1949] <= 16'h6100;
rommem[1950] <= 16'hFFE8;
rommem[1951] <= 16'h6100;
rommem[1952] <= 16'h0092;
rommem[1953] <= 16'h12C1;
rommem[1954] <= 16'h6100;
rommem[1955] <= 16'hFFDE;
rommem[1956] <= 16'h6100;
rommem[1957] <= 16'h0088;
rommem[1958] <= 16'h12C1;
rommem[1959] <= 16'h6100;
rommem[1960] <= 16'hFFD4;
rommem[1961] <= 16'h6100;
rommem[1962] <= 16'h007E;
rommem[1963] <= 16'h12C1;
rommem[1964] <= 16'h6100;
rommem[1965] <= 16'hFFCA;
rommem[1966] <= 16'h6100;
rommem[1967] <= 16'h0074;
rommem[1968] <= 16'h12C1;
rommem[1969] <= 16'h6100;
rommem[1970] <= 16'hFFC0;
rommem[1971] <= 16'h6100;
rommem[1972] <= 16'h006A;
rommem[1973] <= 16'h12C1;
rommem[1974] <= 16'h6100;
rommem[1975] <= 16'hFFB6;
rommem[1976] <= 16'h6100;
rommem[1977] <= 16'h0060;
rommem[1978] <= 16'h12C1;
rommem[1979] <= 16'h6100;
rommem[1980] <= 16'hFFAC;
rommem[1981] <= 16'h6100;
rommem[1982] <= 16'h0056;
rommem[1983] <= 16'h12C1;
rommem[1984] <= 16'h6100;
rommem[1985] <= 16'hFFA2;
rommem[1986] <= 16'h6100;
rommem[1987] <= 16'h004C;
rommem[1988] <= 16'h12C1;
rommem[1989] <= 16'h6000;
rommem[1990] <= 16'hFDF4;
rommem[1991] <= 16'h6100;
rommem[1992] <= 16'hFF94;
rommem[1993] <= 16'h6100;
rommem[1994] <= 16'h003E;
rommem[1995] <= 16'h2041;
rommem[1996] <= 16'h4E90;
rommem[1997] <= 16'h6000;
rommem[1998] <= 16'hFDE4;
rommem[1999] <= 16'h6100;
rommem[2000] <= 16'hFF84;
rommem[2001] <= 16'h6100;
rommem[2002] <= 16'h002E;
rommem[2003] <= 16'h2041;
rommem[2004] <= 16'h4EB9;
rommem[2005] <= 16'hFFFC;
rommem[2006] <= 16'h0232;
rommem[2007] <= 16'h6100;
rommem[2008] <= 16'hF7A2;
rommem[2009] <= 16'h6100;
rommem[2010] <= 16'hF79E;
rommem[2011] <= 16'h6100;
rommem[2012] <= 16'hF79A;
rommem[2013] <= 16'h6100;
rommem[2014] <= 16'hF796;
rommem[2015] <= 16'h6100;
rommem[2016] <= 16'hF792;
rommem[2017] <= 16'h6100;
rommem[2018] <= 16'hF78E;
rommem[2019] <= 16'h6100;
rommem[2020] <= 16'hF78A;
rommem[2021] <= 16'h6100;
rommem[2022] <= 16'hF786;
rommem[2023] <= 16'h6000;
rommem[2024] <= 16'hFDB0;
rommem[2025] <= 16'h48E7;
rommem[2026] <= 16'hA000;
rommem[2027] <= 16'h4282;
rommem[2028] <= 16'h7007;
rommem[2029] <= 16'h1218;
rommem[2030] <= 16'h6100;
rommem[2031] <= 16'h001E;
rommem[2032] <= 16'hB23C;
rommem[2033] <= 16'h00FF;
rommem[2034] <= 16'h670E;
rommem[2035] <= 16'hE98A;
rommem[2036] <= 16'h0281;
rommem[2037] <= 16'h0000;
rommem[2038] <= 16'h000F;
rommem[2039] <= 16'h8481;
rommem[2040] <= 16'h51C8;
rommem[2041] <= 16'hFFE8;
rommem[2042] <= 16'h2202;
rommem[2043] <= 16'h4CDF;
rommem[2044] <= 16'h0005;
rommem[2045] <= 16'h4E75;
rommem[2046] <= 16'h0C01;
rommem[2047] <= 16'h0030;
rommem[2048] <= 16'h6538;
rommem[2049] <= 16'h0C01;
rommem[2050] <= 16'h0039;
rommem[2051] <= 16'h6206;
rommem[2052] <= 16'h0401;
rommem[2053] <= 16'h0030;
rommem[2054] <= 16'h4E75;
rommem[2055] <= 16'h0C01;
rommem[2056] <= 16'h0041;
rommem[2057] <= 16'h6526;
rommem[2058] <= 16'h0C01;
rommem[2059] <= 16'h0046;
rommem[2060] <= 16'h620A;
rommem[2061] <= 16'h0401;
rommem[2062] <= 16'h0041;
rommem[2063] <= 16'h0601;
rommem[2064] <= 16'h000A;
rommem[2065] <= 16'h4E75;
rommem[2066] <= 16'h0C01;
rommem[2067] <= 16'h0061;
rommem[2068] <= 16'h6510;
rommem[2069] <= 16'h0C01;
rommem[2070] <= 16'h0066;
rommem[2071] <= 16'h620A;
rommem[2072] <= 16'h0401;
rommem[2073] <= 16'h0061;
rommem[2074] <= 16'h0601;
rommem[2075] <= 16'h000A;
rommem[2076] <= 16'h4E75;
rommem[2077] <= 16'h72FF;
rommem[2078] <= 16'h4E75;
rommem[2079] <= 16'h4BF9;
rommem[2080] <= 16'hFFE0;
rommem[2081] <= 16'h0000;
rommem[2082] <= 16'h302D;
rommem[2083] <= 16'h04AC;
rommem[2084] <= 16'h0800;
rommem[2085] <= 16'h000D;
rommem[2086] <= 16'h67F6;
rommem[2087] <= 16'h2B7C;
rommem[2088] <= 16'h0001;
rommem[2089] <= 16'hD4C0;
rommem[2090] <= 16'h04BC;
rommem[2091] <= 16'h3B79;
rommem[2092] <= 16'h0001;
rommem[2093] <= 16'h0004;
rommem[2094] <= 16'h04A8;
rommem[2095] <= 16'h2B7C;
rommem[2096] <= 16'h0000;
rommem[2097] <= 16'h0000;
rommem[2098] <= 16'h0498;
rommem[2099] <= 16'h2B7C;
rommem[2100] <= 16'h0000;
rommem[2101] <= 16'h0190;
rommem[2102] <= 16'h04A4;
rommem[2103] <= 16'h2B7C;
rommem[2104] <= 16'h0000;
rommem[2105] <= 16'h0000;
rommem[2106] <= 16'h049C;
rommem[2107] <= 16'h3B7C;
rommem[2108] <= 16'h8080;
rommem[2109] <= 16'h04AC;
rommem[2110] <= 16'h7020;
rommem[2111] <= 16'h323C;
rommem[2112] <= 16'h073A;
rommem[2113] <= 16'h4BF9;
rommem[2114] <= 16'h1FFF;
rommem[2115] <= 16'h0000;
rommem[2116] <= 16'h1AC0;
rommem[2117] <= 16'h51C9;
rommem[2118] <= 16'hFFFC;
rommem[2119] <= 16'h4E75;
rommem[2120] <= 16'h48E7;
rommem[2121] <= 16'h8084;
rommem[2122] <= 16'h4BF9;
rommem[2123] <= 16'hFFE0;
rommem[2124] <= 16'h0000;
rommem[2125] <= 16'h302D;
rommem[2126] <= 16'h04AC;
rommem[2127] <= 16'h0800;
rommem[2128] <= 16'h000D;
rommem[2129] <= 16'h67F6;
rommem[2130] <= 16'h2B7C;
rommem[2131] <= 16'h0001;
rommem[2132] <= 16'hC840;
rommem[2133] <= 16'h04B0;
rommem[2134] <= 16'h2B7C;
rommem[2135] <= 16'h0000;
rommem[2136] <= 16'h0C80;
rommem[2137] <= 16'h0480;
rommem[2138] <= 16'h2B7C;
rommem[2139] <= 16'h0000;
rommem[2140] <= 16'h0000;
rommem[2141] <= 16'h0484;
rommem[2142] <= 16'h2B7C;
rommem[2143] <= 16'h0001;
rommem[2144] <= 16'hC840;
rommem[2145] <= 16'h04BC;
rommem[2146] <= 16'h2B7C;
rommem[2147] <= 16'h0000;
rommem[2148] <= 16'h0000;
rommem[2149] <= 16'h0498;
rommem[2150] <= 16'h2B7C;
rommem[2151] <= 16'h0000;
rommem[2152] <= 16'h0000;
rommem[2153] <= 16'h049C;
rommem[2154] <= 16'h2B7C;
rommem[2155] <= 16'hFFFF;
rommem[2156] <= 16'hFFFF;
rommem[2157] <= 16'h04A0;
rommem[2158] <= 16'h2B7C;
rommem[2159] <= 16'hFFFF;
rommem[2160] <= 16'hFFFF;
rommem[2161] <= 16'h04A4;
rommem[2162] <= 16'h3B7C;
rommem[2163] <= 16'h0011;
rommem[2164] <= 16'h04AE;
rommem[2165] <= 16'h3B7C;
rommem[2166] <= 16'h8082;
rommem[2167] <= 16'h04AC;
rommem[2168] <= 16'h4BF9;
rommem[2169] <= 16'h1FFF;
rommem[2170] <= 16'h0000;
rommem[2171] <= 16'h204D;
rommem[2172] <= 16'h1039;
rommem[2173] <= 16'h0001;
rommem[2174] <= 16'h041B;
rommem[2175] <= 16'h4880;
rommem[2176] <= 16'hD1C0;
rommem[2177] <= 16'hC0FC;
rommem[2178] <= 16'h0025;
rommem[2179] <= 16'h1AD8;
rommem[2180] <= 16'h51C8;
rommem[2181] <= 16'hFFFC;
rommem[2182] <= 16'h4CDF;
rommem[2183] <= 16'h2101;
rommem[2184] <= 16'h48E7;
rommem[2185] <= 16'h8004;
rommem[2186] <= 16'h4BF9;
rommem[2187] <= 16'hFFE0;
rommem[2188] <= 16'h0000;
rommem[2189] <= 16'h302D;
rommem[2190] <= 16'h04AC;
rommem[2191] <= 16'h0800;
rommem[2192] <= 16'h000D;
rommem[2193] <= 16'h67F6;
rommem[2194] <= 16'h2B7C;
rommem[2195] <= 16'h0000;
rommem[2196] <= 16'h0C80;
rommem[2197] <= 16'h04BC;
rommem[2198] <= 16'h2B7C;
rommem[2199] <= 16'h0001;
rommem[2200] <= 16'hC840;
rommem[2201] <= 16'h0498;
rommem[2202] <= 16'h2B7C;
rommem[2203] <= 16'h0000;
rommem[2204] <= 16'h0000;
rommem[2205] <= 16'h049C;
rommem[2206] <= 16'h2B7C;
rommem[2207] <= 16'hFFFF;
rommem[2208] <= 16'hFFFF;
rommem[2209] <= 16'h04A4;
rommem[2210] <= 16'h3B79;
rommem[2211] <= 16'h0001;
rommem[2212] <= 16'h0004;
rommem[2213] <= 16'h04A8;
rommem[2214] <= 16'h3B7C;
rommem[2215] <= 16'h8080;
rommem[2216] <= 16'h04AC;
rommem[2217] <= 16'h4BF9;
rommem[2218] <= 16'h1FFF;
rommem[2219] <= 16'h073A;
rommem[2220] <= 16'h7028;
rommem[2221] <= 16'h1AFC;
rommem[2222] <= 16'h0020;
rommem[2223] <= 16'h51C8;
rommem[2224] <= 16'hFFFA;
rommem[2225] <= 16'h4CDF;
rommem[2226] <= 16'h2001;
rommem[2227] <= 16'h4E75;
rommem[2228] <= 16'h600A;
rommem[2229] <= 16'h6100;
rommem[2230] <= 16'h017A;
rommem[2231] <= 16'h0C00;
rommem[2232] <= 16'h000A;
rommem[2233] <= 16'h66F6;
rommem[2234] <= 16'h6100;
rommem[2235] <= 16'h0170;
rommem[2236] <= 16'h1800;
rommem[2237] <= 16'h0C04;
rommem[2238] <= 16'h001A;
rommem[2239] <= 16'h6700;
rommem[2240] <= 16'hFC00;
rommem[2241] <= 16'h0C04;
rommem[2242] <= 16'h0053;
rommem[2243] <= 16'h66E2;
rommem[2244] <= 16'h6100;
rommem[2245] <= 16'h015C;
rommem[2246] <= 16'h1800;
rommem[2247] <= 16'h0C04;
rommem[2248] <= 16'h0030;
rommem[2249] <= 16'h65D6;
rommem[2250] <= 16'h0C04;
rommem[2251] <= 16'h0039;
rommem[2252] <= 16'h62D0;
rommem[2253] <= 16'h6100;
rommem[2254] <= 16'h014A;
rommem[2255] <= 16'h6100;
rommem[2256] <= 16'hFE5C;
rommem[2257] <= 16'h1401;
rommem[2258] <= 16'h6100;
rommem[2259] <= 16'h0140;
rommem[2260] <= 16'h6100;
rommem[2261] <= 16'hFE52;
rommem[2262] <= 16'hE90A;
rommem[2263] <= 16'h8202;
rommem[2264] <= 16'h1601;
rommem[2265] <= 16'h0C04;
rommem[2266] <= 16'h0030;
rommem[2267] <= 16'h67B2;
rommem[2268] <= 16'h0C04;
rommem[2269] <= 16'h0031;
rommem[2270] <= 16'h676A;
rommem[2271] <= 16'h0C04;
rommem[2272] <= 16'h0032;
rommem[2273] <= 16'h676A;
rommem[2274] <= 16'h0C04;
rommem[2275] <= 16'h0033;
rommem[2276] <= 16'h676A;
rommem[2277] <= 16'h0C04;
rommem[2278] <= 16'h0035;
rommem[2279] <= 16'h679A;
rommem[2280] <= 16'h0C04;
rommem[2281] <= 16'h0037;
rommem[2282] <= 16'h6764;
rommem[2283] <= 16'h0C04;
rommem[2284] <= 16'h0038;
rommem[2285] <= 16'h676C;
rommem[2286] <= 16'h0C04;
rommem[2287] <= 16'h0039;
rommem[2288] <= 16'h6774;
rommem[2289] <= 16'h6086;
rommem[2290] <= 16'h0243;
rommem[2291] <= 16'h00FF;
rommem[2292] <= 16'h5343;
rommem[2293] <= 16'h4282;
rommem[2294] <= 16'h6100;
rommem[2295] <= 16'h00F8;
rommem[2296] <= 16'h6100;
rommem[2297] <= 16'hFE0A;
rommem[2298] <= 16'hE98A;
rommem[2299] <= 16'h8401;
rommem[2300] <= 16'h6100;
rommem[2301] <= 16'h00EC;
rommem[2302] <= 16'h6100;
rommem[2303] <= 16'hFDFE;
rommem[2304] <= 16'hE98A;
rommem[2305] <= 16'h8401;
rommem[2306] <= 16'h12C2;
rommem[2307] <= 16'h51CB;
rommem[2308] <= 16'hFFE2;
rommem[2309] <= 16'h4282;
rommem[2310] <= 16'h6100;
rommem[2311] <= 16'h00D8;
rommem[2312] <= 16'h6100;
rommem[2313] <= 16'hFDEA;
rommem[2314] <= 16'hE98A;
rommem[2315] <= 16'h8401;
rommem[2316] <= 16'h6100;
rommem[2317] <= 16'h00CC;
rommem[2318] <= 16'h6100;
rommem[2319] <= 16'hFDDE;
rommem[2320] <= 16'hE98A;
rommem[2321] <= 16'h8401;
rommem[2322] <= 16'h6000;
rommem[2323] <= 16'hFF44;
rommem[2324] <= 16'h6100;
rommem[2325] <= 16'h003A;
rommem[2326] <= 16'h60B6;
rommem[2327] <= 16'h6100;
rommem[2328] <= 16'h0042;
rommem[2329] <= 16'h60B0;
rommem[2330] <= 16'h6100;
rommem[2331] <= 16'h004A;
rommem[2332] <= 16'h60AA;
rommem[2333] <= 16'h6100;
rommem[2334] <= 16'h0044;
rommem[2335] <= 16'h23C9;
rommem[2336] <= 16'h0000;
rommem[2337] <= 16'h0000;
rommem[2338] <= 16'h6000;
rommem[2339] <= 16'hFB3A;
rommem[2340] <= 16'h6100;
rommem[2341] <= 16'h0028;
rommem[2342] <= 16'h23C9;
rommem[2343] <= 16'h0000;
rommem[2344] <= 16'h0000;
rommem[2345] <= 16'h6000;
rommem[2346] <= 16'hFB2C;
rommem[2347] <= 16'h6100;
rommem[2348] <= 16'h000C;
rommem[2349] <= 16'h23C9;
rommem[2350] <= 16'h0000;
rommem[2351] <= 16'h0000;
rommem[2352] <= 16'h6000;
rommem[2353] <= 16'hFB1E;
rommem[2354] <= 16'h4282;
rommem[2355] <= 16'h6100;
rommem[2356] <= 16'h007E;
rommem[2357] <= 16'h6100;
rommem[2358] <= 16'hFD90;
rommem[2359] <= 16'h1401;
rommem[2360] <= 16'h604A;
rommem[2361] <= 16'h4282;
rommem[2362] <= 16'h6100;
rommem[2363] <= 16'h0070;
rommem[2364] <= 16'h6100;
rommem[2365] <= 16'hFD82;
rommem[2366] <= 16'h1401;
rommem[2367] <= 16'h6024;
rommem[2368] <= 16'h4282;
rommem[2369] <= 16'h6100;
rommem[2370] <= 16'h0062;
rommem[2371] <= 16'h6100;
rommem[2372] <= 16'hFD74;
rommem[2373] <= 16'h1401;
rommem[2374] <= 16'h6100;
rommem[2375] <= 16'h0058;
rommem[2376] <= 16'h6100;
rommem[2377] <= 16'hFD6A;
rommem[2378] <= 16'hE98A;
rommem[2379] <= 16'h8401;
rommem[2380] <= 16'h6100;
rommem[2381] <= 16'h004C;
rommem[2382] <= 16'h6100;
rommem[2383] <= 16'hFD5E;
rommem[2384] <= 16'hE98A;
rommem[2385] <= 16'h8401;
rommem[2386] <= 16'h6100;
rommem[2387] <= 16'h0040;
rommem[2388] <= 16'h6100;
rommem[2389] <= 16'hFD52;
rommem[2390] <= 16'hE98A;
rommem[2391] <= 16'h8401;
rommem[2392] <= 16'h6100;
rommem[2393] <= 16'h0034;
rommem[2394] <= 16'h6100;
rommem[2395] <= 16'hFD46;
rommem[2396] <= 16'hE98A;
rommem[2397] <= 16'h8401;
rommem[2398] <= 16'h6100;
rommem[2399] <= 16'h0028;
rommem[2400] <= 16'h6100;
rommem[2401] <= 16'hFD3A;
rommem[2402] <= 16'hE98A;
rommem[2403] <= 16'h8401;
rommem[2404] <= 16'h6100;
rommem[2405] <= 16'h001C;
rommem[2406] <= 16'h6100;
rommem[2407] <= 16'hFD2E;
rommem[2408] <= 16'hE98A;
rommem[2409] <= 16'h8401;
rommem[2410] <= 16'h6100;
rommem[2411] <= 16'h0010;
rommem[2412] <= 16'h6100;
rommem[2413] <= 16'hFD22;
rommem[2414] <= 16'hE98A;
rommem[2415] <= 16'h8401;
rommem[2416] <= 16'h4284;
rommem[2417] <= 16'h2242;
rommem[2418] <= 16'h4E75;
rommem[2419] <= 16'h6100;
rommem[2420] <= 16'hF500;
rommem[2421] <= 16'h670C;
rommem[2422] <= 16'h6100;
rommem[2423] <= 16'hF50C;
rommem[2424] <= 16'h0C01;
rommem[2425] <= 16'h0003;
rommem[2426] <= 16'h6700;
rommem[2427] <= 16'hFA8A;
rommem[2428] <= 16'h6100;
rommem[2429] <= 16'hFFFF;
rommem[2430] <= 16'h67E8;
rommem[2431] <= 16'h1200;
rommem[2432] <= 16'h4E75;
rommem[2433] <= 16'h33FC;
rommem[2434] <= 16'hA6A6;
rommem[2435] <= 16'hFFDC;
rommem[2436] <= 16'h0600;
rommem[2437] <= 16'h2C7C;
rommem[2438] <= 16'hFFE0;
rommem[2439] <= 16'h0000;
rommem[2440] <= 16'h343C;
rommem[2441] <= 16'h0007;
rommem[2442] <= 16'h1001;
rommem[2443] <= 16'h0240;
rommem[2444] <= 16'h000F;
rommem[2445] <= 16'h0C40;
rommem[2446] <= 16'h0009;
rommem[2447] <= 16'h6302;
rommem[2448] <= 16'h5E40;
rommem[2449] <= 16'h0640;
rommem[2450] <= 16'h0030;
rommem[2451] <= 16'h3602;
rommem[2452] <= 16'hE743;
rommem[2453] <= 16'h382E;
rommem[2454] <= 16'h042C;
rommem[2455] <= 16'hB87C;
rommem[2456] <= 16'h001C;
rommem[2457] <= 16'h64F6;
rommem[2458] <= 16'h4880;
rommem[2459] <= 16'h3D40;
rommem[2460] <= 16'h0420;
rommem[2461] <= 16'h3D7C;
rommem[2462] <= 16'h7FFF;
rommem[2463] <= 16'h0422;
rommem[2464] <= 16'h3D7C;
rommem[2465] <= 16'h000F;
rommem[2466] <= 16'h0424;
rommem[2467] <= 16'h3D43;
rommem[2468] <= 16'h0426;
rommem[2469] <= 16'h3D7C;
rommem[2470] <= 16'h0008;
rommem[2471] <= 16'h0428;
rommem[2472] <= 16'h3D7C;
rommem[2473] <= 16'h0707;
rommem[2474] <= 16'h042A;
rommem[2475] <= 16'h3D7C;
rommem[2476] <= 16'h0000;
rommem[2477] <= 16'h042E;
rommem[2478] <= 16'hE899;
rommem[2479] <= 16'h57CA;
rommem[2480] <= 16'hFFB4;
rommem[2481] <= 16'h4ED5;
rommem[2482] <= 16'h33FC;
rommem[2483] <= 16'hA5A5;
rommem[2484] <= 16'hFFDC;
rommem[2485] <= 16'h0600;
rommem[2486] <= 16'h207C;
rommem[2487] <= 16'h0003;
rommem[2488] <= 16'h0000;
rommem[2489] <= 16'h203C;
rommem[2490] <= 16'hAAAA;
rommem[2491] <= 16'h5555;
rommem[2492] <= 16'h20C0;
rommem[2493] <= 16'h2208;
rommem[2494] <= 16'h4A41;
rommem[2495] <= 16'h660A;
rommem[2496] <= 16'h4BF9;
rommem[2497] <= 16'hFFFC;
rommem[2498] <= 16'h138A;
rommem[2499] <= 16'h6000;
rommem[2500] <= 16'hFF7A;
rommem[2501] <= 16'h33FC;
rommem[2502] <= 16'hA9A9;
rommem[2503] <= 16'hFFDC;
rommem[2504] <= 16'h0600;
rommem[2505] <= 16'hB1FC;
rommem[2506] <= 16'h0005;
rommem[2507] <= 16'hFFFC;
rommem[2508] <= 16'h66DE;
rommem[2509] <= 16'h7200;
rommem[2510] <= 16'h6100;
rommem[2511] <= 16'hEEAE;
rommem[2512] <= 16'h6000;
rommem[2513] <= 16'hFC04;
rommem[2514] <= 16'h33FC;
rommem[2515] <= 16'hA7A7;
rommem[2516] <= 16'hFFDC;
rommem[2517] <= 16'h0600;
rommem[2518] <= 16'h2448;
rommem[2519] <= 16'h207C;
rommem[2520] <= 16'h0003;
rommem[2521] <= 16'h0000;
rommem[2522] <= 16'h2A18;
rommem[2523] <= 16'hB5C8;
rommem[2524] <= 16'h671A;
rommem[2525] <= 16'h2208;
rommem[2526] <= 16'h4A41;
rommem[2527] <= 16'h660A;
rommem[2528] <= 16'h4BF9;
rommem[2529] <= 16'hFFFC;
rommem[2530] <= 16'h13CA;
rommem[2531] <= 16'h6000;
rommem[2532] <= 16'hFF3A;
rommem[2533] <= 16'h0C85;
rommem[2534] <= 16'hAAAA;
rommem[2535] <= 16'h5555;
rommem[2536] <= 16'h67E2;
rommem[2537] <= 16'h6678;
rommem[2538] <= 16'h33FC;
rommem[2539] <= 16'hA8A8;
rommem[2540] <= 16'hFFDC;
rommem[2541] <= 16'h0600;
rommem[2542] <= 16'h207C;
rommem[2543] <= 16'h0003;
rommem[2544] <= 16'h0000;
rommem[2545] <= 16'h203C;
rommem[2546] <= 16'h5555;
rommem[2547] <= 16'hAAAA;
rommem[2548] <= 16'h20C0;
rommem[2549] <= 16'h2208;
rommem[2550] <= 16'h4A41;
rommem[2551] <= 16'h660A;
rommem[2552] <= 16'h4BF9;
rommem[2553] <= 16'hFFFC;
rommem[2554] <= 16'h13FA;
rommem[2555] <= 16'h6000;
rommem[2556] <= 16'hFF0A;
rommem[2557] <= 16'hB1FC;
rommem[2558] <= 16'h1FFF;
rommem[2559] <= 16'hFFFC;
rommem[2560] <= 16'h66E6;
rommem[2561] <= 16'h2448;
rommem[2562] <= 16'h207C;
rommem[2563] <= 16'h0003;
rommem[2564] <= 16'h0000;
rommem[2565] <= 16'h2018;
rommem[2566] <= 16'hB5C8;
rommem[2567] <= 16'h671A;
rommem[2568] <= 16'h2208;
rommem[2569] <= 16'h4A41;
rommem[2570] <= 16'h660A;
rommem[2571] <= 16'h4BF9;
rommem[2572] <= 16'hFFFC;
rommem[2573] <= 16'h1420;
rommem[2574] <= 16'h6000;
rommem[2575] <= 16'hFEE4;
rommem[2576] <= 16'h0C80;
rommem[2577] <= 16'h5555;
rommem[2578] <= 16'hAAAA;
rommem[2579] <= 16'h67E2;
rommem[2580] <= 16'h6622;
rommem[2581] <= 16'h23C8;
rommem[2582] <= 16'h0001;
rommem[2583] <= 16'h0008;
rommem[2584] <= 16'h91FC;
rommem[2585] <= 16'h0000;
rommem[2586] <= 16'h000C;
rommem[2587] <= 16'h21C8;
rommem[2588] <= 16'h0404;
rommem[2589] <= 16'h21FC;
rommem[2590] <= 16'h4652;
rommem[2591] <= 16'h4545;
rommem[2592] <= 16'h0400;
rommem[2593] <= 16'h21FC;
rommem[2594] <= 16'h0000;
rommem[2595] <= 16'h0408;
rommem[2596] <= 16'h0408;
rommem[2597] <= 16'h4ED3;
rommem[2598] <= 16'h4ED3;
rommem[2599] <= 16'h60FC;
rommem[2600] <= 16'h6100;
rommem[2601] <= 16'h0080;
rommem[2602] <= 16'h6100;
rommem[2603] <= 16'h0006;
rommem[2604] <= 16'h6000;
rommem[2605] <= 16'hF926;
rommem[2606] <= 16'h4DF9;
rommem[2607] <= 16'hFFDC;
rommem[2608] <= 16'h0000;
rommem[2609] <= 16'h4BF9;
rommem[2610] <= 16'hFFE0;
rommem[2611] <= 16'h0000;
rommem[2612] <= 16'h2C3C;
rommem[2613] <= 16'h0000;
rommem[2614] <= 16'h4E20;
rommem[2615] <= 16'h202E;
rommem[2616] <= 16'h0C00;
rommem[2617] <= 16'h3200;
rommem[2618] <= 16'h4840;
rommem[2619] <= 16'h0240;
rommem[2620] <= 16'h00FF;
rommem[2621] <= 16'h0241;
rommem[2622] <= 16'h00FF;
rommem[2623] <= 16'h426E;
rommem[2624] <= 16'h0C04;
rommem[2625] <= 16'h242E;
rommem[2626] <= 16'h0C00;
rommem[2627] <= 16'h3602;
rommem[2628] <= 16'h4842;
rommem[2629] <= 16'h0242;
rommem[2630] <= 16'h00FF;
rommem[2631] <= 16'h0243;
rommem[2632] <= 16'h00FF;
rommem[2633] <= 16'h426E;
rommem[2634] <= 16'h0C04;
rommem[2635] <= 16'h282E;
rommem[2636] <= 16'h0C00;
rommem[2637] <= 16'h0244;
rommem[2638] <= 16'h7FFF;
rommem[2639] <= 16'h426E;
rommem[2640] <= 16'h0C04;
rommem[2641] <= 16'h3E2D;
rommem[2642] <= 16'h042C;
rommem[2643] <= 16'hBE7C;
rommem[2644] <= 16'h001C;
rommem[2645] <= 16'h64F6;
rommem[2646] <= 16'h3B7C;
rommem[2647] <= 16'h0001;
rommem[2648] <= 16'h0422;
rommem[2649] <= 16'h3B44;
rommem[2650] <= 16'h0424;
rommem[2651] <= 16'h3B40;
rommem[2652] <= 16'h0426;
rommem[2653] <= 16'h3B41;
rommem[2654] <= 16'h0428;
rommem[2655] <= 16'h3B42;
rommem[2656] <= 16'h0430;
rommem[2657] <= 16'h3B43;
rommem[2658] <= 16'h0432;
rommem[2659] <= 16'h3B7C;
rommem[2660] <= 16'h0003;
rommem[2661] <= 16'h042E;
rommem[2662] <= 16'h5386;
rommem[2663] <= 16'h669E;
rommem[2664] <= 16'h4E75;
rommem[2665] <= 16'h4DF9;
rommem[2666] <= 16'hFFDC;
rommem[2667] <= 16'h0000;
rommem[2668] <= 16'h4BF9;
rommem[2669] <= 16'hFFE0;
rommem[2670] <= 16'h0000;
rommem[2671] <= 16'h2C3C;
rommem[2672] <= 16'h0003;
rommem[2673] <= 16'h0D40;
rommem[2674] <= 16'h33FC;
rommem[2675] <= 16'h000A;
rommem[2676] <= 16'hFFDC;
rommem[2677] <= 16'h0600;
rommem[2678] <= 16'h302D;
rommem[2679] <= 16'h04AC;
rommem[2680] <= 16'h0800;
rommem[2681] <= 16'h000E;
rommem[2682] <= 16'h6706;
rommem[2683] <= 16'h0800;
rommem[2684] <= 16'h000D;
rommem[2685] <= 16'h67E8;
rommem[2686] <= 16'h33FC;
rommem[2687] <= 16'h000B;
rommem[2688] <= 16'hFFDC;
rommem[2689] <= 16'h0600;
rommem[2690] <= 16'h202E;
rommem[2691] <= 16'h0C00;
rommem[2692] <= 16'h3200;
rommem[2693] <= 16'h4840;
rommem[2694] <= 16'h0240;
rommem[2695] <= 16'h00FF;
rommem[2696] <= 16'h0241;
rommem[2697] <= 16'h00FF;
rommem[2698] <= 16'h426E;
rommem[2699] <= 16'h0C04;
rommem[2700] <= 16'h242E;
rommem[2701] <= 16'h0C00;
rommem[2702] <= 16'h3602;
rommem[2703] <= 16'h4842;
rommem[2704] <= 16'h0242;
rommem[2705] <= 16'h00FF;
rommem[2706] <= 16'h0243;
rommem[2707] <= 16'h00FF;
rommem[2708] <= 16'h426E;
rommem[2709] <= 16'h0C04;
rommem[2710] <= 16'h282E;
rommem[2711] <= 16'h0C00;
rommem[2712] <= 16'h0244;
rommem[2713] <= 16'h7FFF;
rommem[2714] <= 16'h426E;
rommem[2715] <= 16'h0C04;
rommem[2716] <= 16'h3E2D;
rommem[2717] <= 16'h042C;
rommem[2718] <= 16'hBE7C;
rommem[2719] <= 16'h001C;
rommem[2720] <= 16'h64F6;
rommem[2721] <= 16'h33FC;
rommem[2722] <= 16'h000C;
rommem[2723] <= 16'hFFDC;
rommem[2724] <= 16'h0600;
rommem[2725] <= 16'h3B7C;
rommem[2726] <= 16'h0001;
rommem[2727] <= 16'h0422;
rommem[2728] <= 16'h3B44;
rommem[2729] <= 16'h0424;
rommem[2730] <= 16'h3B40;
rommem[2731] <= 16'h0426;
rommem[2732] <= 16'h3B41;
rommem[2733] <= 16'h0428;
rommem[2734] <= 16'h3B42;
rommem[2735] <= 16'h0430;
rommem[2736] <= 16'h3B43;
rommem[2737] <= 16'h0432;
rommem[2738] <= 16'h3B7C;
rommem[2739] <= 16'h0002;
rommem[2740] <= 16'h042E;
rommem[2741] <= 16'h5386;
rommem[2742] <= 16'h6600;
rommem[2743] <= 16'hFF76;
rommem[2744] <= 16'h4E75;
rommem[2745] <= 16'h4BF9;
rommem[2746] <= 16'hFFE0;
rommem[2747] <= 16'h0000;
rommem[2748] <= 16'h302D;
rommem[2749] <= 16'h04AC;
rommem[2750] <= 16'h0800;
rommem[2751] <= 16'h000D;
rommem[2752] <= 16'h67F6;
rommem[2753] <= 16'h2B7C;
rommem[2754] <= 16'h0000;
rommem[2755] <= 16'h1F40;
rommem[2756] <= 16'h04BC;
rommem[2757] <= 16'h3B7C;
rommem[2758] <= 16'h7C00;
rommem[2759] <= 16'h04A8;
rommem[2760] <= 16'h2B7C;
rommem[2761] <= 16'h0000;
rommem[2762] <= 16'h0168;
rommem[2763] <= 16'h0498;
rommem[2764] <= 16'h2B7C;
rommem[2765] <= 16'h0000;
rommem[2766] <= 16'h0028;
rommem[2767] <= 16'h04A4;
rommem[2768] <= 16'h2B7C;
rommem[2769] <= 16'h0000;
rommem[2770] <= 16'h0168;
rommem[2771] <= 16'h049C;
rommem[2772] <= 16'h3B7C;
rommem[2773] <= 16'h8080;
rommem[2774] <= 16'h04AC;
rommem[2775] <= 16'h302D;
rommem[2776] <= 16'h04AC;
rommem[2777] <= 16'h0800;
rommem[2778] <= 16'h000D;
rommem[2779] <= 16'h67F6;
rommem[2780] <= 16'h2B7C;
rommem[2781] <= 16'h0000;
rommem[2782] <= 16'h03E8;
rommem[2783] <= 16'h04B0;
rommem[2784] <= 16'h2B7C;
rommem[2785] <= 16'h0000;
rommem[2786] <= 16'h0000;
rommem[2787] <= 16'h0480;
rommem[2788] <= 16'h2B7C;
rommem[2789] <= 16'h0000;
rommem[2790] <= 16'h0168;
rommem[2791] <= 16'h0484;
rommem[2792] <= 16'h2B7C;
rommem[2793] <= 16'h0000;
rommem[2794] <= 16'h03E8;
rommem[2795] <= 16'h04B8;
rommem[2796] <= 16'h2B7C;
rommem[2797] <= 16'h0000;
rommem[2798] <= 16'h0000;
rommem[2799] <= 16'h0490;
rommem[2800] <= 16'h2B7C;
rommem[2801] <= 16'h0000;
rommem[2802] <= 16'h0168;
rommem[2803] <= 16'h0494;
rommem[2804] <= 16'h2B7C;
rommem[2805] <= 16'h0000;
rommem[2806] <= 16'h1F40;
rommem[2807] <= 16'h04BC;
rommem[2808] <= 16'h2B7C;
rommem[2809] <= 16'h0000;
rommem[2810] <= 16'h0140;
rommem[2811] <= 16'h0498;
rommem[2812] <= 16'h2B7C;
rommem[2813] <= 16'h0000;
rommem[2814] <= 16'h0168;
rommem[2815] <= 16'h049C;
rommem[2816] <= 16'h2B7C;
rommem[2817] <= 16'h0000;
rommem[2818] <= 16'h0028;
rommem[2819] <= 16'h04A0;
rommem[2820] <= 16'h2B7C;
rommem[2821] <= 16'h0000;
rommem[2822] <= 16'h0028;
rommem[2823] <= 16'h04A4;
rommem[2824] <= 16'h3B7C;
rommem[2825] <= 16'h0091;
rommem[2826] <= 16'h04AE;
rommem[2827] <= 16'h3B7C;
rommem[2828] <= 16'h80A2;
rommem[2829] <= 16'h04AC;
rommem[2830] <= 16'h302D;
rommem[2831] <= 16'h04AC;
rommem[2832] <= 16'h0800;
rommem[2833] <= 16'h000D;
rommem[2834] <= 16'h67F6;
rommem[2835] <= 16'h4E75;
rommem[2836] <= 16'h4DF9;
rommem[2837] <= 16'hFFDC;
rommem[2838] <= 16'h0E00;
rommem[2839] <= 16'h3CBC;
rommem[2840] <= 16'h0013;
rommem[2841] <= 16'h3D7C;
rommem[2842] <= 16'h0000;
rommem[2843] <= 16'h0002;
rommem[2844] <= 16'h4DF9;
rommem[2845] <= 16'hFFDC;
rommem[2846] <= 16'h0E10;
rommem[2847] <= 16'h3CBC;
rommem[2848] <= 16'h0013;
rommem[2849] <= 16'h3D7C;
rommem[2850] <= 16'h0000;
rommem[2851] <= 16'h0002;
rommem[2852] <= 16'h4E75;
rommem[2853] <= 16'h3F00;
rommem[2854] <= 16'h302E;
rommem[2855] <= 16'h000A;
rommem[2856] <= 16'h0800;
rommem[2857] <= 16'h0001;
rommem[2858] <= 16'h66F6;
rommem[2859] <= 16'h301F;
rommem[2860] <= 16'h4E75;
rommem[2861] <= 16'h3D40;
rommem[2862] <= 16'h0006;
rommem[2863] <= 16'h3D41;
rommem[2864] <= 16'h0008;
rommem[2865] <= 16'h6100;
rommem[2866] <= 16'hFFE6;
rommem[2867] <= 16'h302E;
rommem[2868] <= 16'h000A;
rommem[2869] <= 16'h4E75;
rommem[2870] <= 16'h3F00;
rommem[2871] <= 16'h3D7C;
rommem[2872] <= 16'h0001;
rommem[2873] <= 16'h0004;
rommem[2874] <= 16'h7076;
rommem[2875] <= 16'h323C;
rommem[2876] <= 16'h0090;
rommem[2877] <= 16'h6100;
rommem[2878] <= 16'hFFDE;
rommem[2879] <= 16'h6100;
rommem[2880] <= 16'h0010;
rommem[2881] <= 16'h301F;
rommem[2882] <= 16'h323C;
rommem[2883] <= 16'h0050;
rommem[2884] <= 16'h6100;
rommem[2885] <= 16'hFFD0;
rommem[2886] <= 16'h6100;
rommem[2887] <= 16'h0002;
rommem[2888] <= 16'h3F00;
rommem[2889] <= 16'h302E;
rommem[2890] <= 16'h000A;
rommem[2891] <= 16'h0800;
rommem[2892] <= 16'h0007;
rommem[2893] <= 16'h66F6;
rommem[2894] <= 16'h301F;
rommem[2895] <= 16'h4E75;
rommem[2896] <= 16'h4BF9;
rommem[2897] <= 16'hFFE0;
rommem[2898] <= 16'h0000;
rommem[2899] <= 16'h2B7C;
rommem[2900] <= 16'h0005;
rommem[2901] <= 16'h8000;
rommem[2902] <= 16'h0640;
rommem[2903] <= 16'h3B7C;
rommem[2904] <= 16'h4000;
rommem[2905] <= 16'h0644;
rommem[2906] <= 16'h3B7C;
rommem[2907] <= 16'h0716;
rommem[2908] <= 16'h0646;
rommem[2909] <= 16'h3B7C;
rommem[2910] <= 16'h1090;
rommem[2911] <= 16'h0584;
rommem[2912] <= 16'h3B7C;
rommem[2913] <= 16'h0090;
rommem[2914] <= 16'h0584;
rommem[2915] <= 16'h302D;
rommem[2916] <= 16'h04AC;
rommem[2917] <= 16'h0800;
rommem[2918] <= 16'h000D;
rommem[2919] <= 16'h67F6;
rommem[2920] <= 16'h2B7C;
rommem[2921] <= 16'h0001;
rommem[2922] <= 16'h0000;
rommem[2923] <= 16'h04BC;
rommem[2924] <= 16'h3B7C;
rommem[2925] <= 16'h000F;
rommem[2926] <= 16'h04A8;
rommem[2927] <= 16'h2B7C;
rommem[2928] <= 16'h0000;
rommem[2929] <= 16'h0000;
rommem[2930] <= 16'h0498;
rommem[2931] <= 16'h2B7C;
rommem[2932] <= 16'h0000;
rommem[2933] <= 16'h0100;
rommem[2934] <= 16'h04A4;
rommem[2935] <= 16'h2B7C;
rommem[2936] <= 16'h0000;
rommem[2937] <= 16'h0040;
rommem[2938] <= 16'h049C;
rommem[2939] <= 16'h3B7C;
rommem[2940] <= 16'h8080;
rommem[2941] <= 16'h04AC;
rommem[2942] <= 16'h203C;
rommem[2943] <= 16'h0003;
rommem[2944] <= 16'hD090;
rommem[2945] <= 16'h5380;
rommem[2946] <= 16'h66FC;
rommem[2947] <= 16'h60BE;
rommem[2948] <= 16'h7000;
rommem[2949] <= 16'h720E;
rommem[2950] <= 16'h6100;
rommem[2951] <= 16'h001C;
rommem[2952] <= 16'h7002;
rommem[2953] <= 16'h41F9;
rommem[2954] <= 16'hFFFC;
rommem[2955] <= 16'h1784;
rommem[2956] <= 16'h6100;
rommem[2957] <= 16'h0076;
rommem[2958] <= 16'h4E75;
rommem[2959] <= 16'h4E75;
rommem[2960] <= 16'h6100;
rommem[2961] <= 16'hFFE6;
rommem[2962] <= 16'h6100;
rommem[2963] <= 16'hFFF8;
rommem[2964] <= 16'h4E75;
rommem[2965] <= 16'h4DF9;
rommem[2966] <= 16'hFFDC;
rommem[2967] <= 16'h0E00;
rommem[2968] <= 16'h3D7C;
rommem[2969] <= 16'h0001;
rommem[2970] <= 16'h0004;
rommem[2971] <= 16'h3D7C;
rommem[2972] <= 16'h0076;
rommem[2973] <= 16'h0006;
rommem[2974] <= 16'h3D7C;
rommem[2975] <= 16'h0090;
rommem[2976] <= 16'h0008;
rommem[2977] <= 16'h6100;
rommem[2978] <= 16'hFF06;
rommem[2979] <= 16'h6100;
rommem[2980] <= 16'hFF48;
rommem[2981] <= 16'h3D7C;
rommem[2982] <= 16'h0040;
rommem[2983] <= 16'h0006;
rommem[2984] <= 16'h3D7C;
rommem[2985] <= 16'h0010;
rommem[2986] <= 16'h0008;
rommem[2987] <= 16'h6100;
rommem[2988] <= 16'hFEF2;
rommem[2989] <= 16'h6100;
rommem[2990] <= 16'hFF34;
rommem[2991] <= 16'h3D40;
rommem[2992] <= 16'h0006;
rommem[2993] <= 16'h3D7C;
rommem[2994] <= 16'h0010;
rommem[2995] <= 16'h0008;
rommem[2996] <= 16'h6100;
rommem[2997] <= 16'hFEE0;
rommem[2998] <= 16'h6100;
rommem[2999] <= 16'hFF22;
rommem[3000] <= 16'h3D41;
rommem[3001] <= 16'h0006;
rommem[3002] <= 16'h3D7C;
rommem[3003] <= 16'h0050;
rommem[3004] <= 16'h0008;
rommem[3005] <= 16'h6100;
rommem[3006] <= 16'hFECE;
rommem[3007] <= 16'h6100;
rommem[3008] <= 16'hFF10;
rommem[3009] <= 16'h4E75;
rommem[3010] <= 16'h0000;
rommem[3011] <= 16'h007D;
rommem[3012] <= 16'h0000;
rommem[3013] <= 16'h000C;
rommem[3014] <= 16'h0020;
rommem[3015] <= 16'h0001;
rommem[3016] <= 16'h41F9;
rommem[3017] <= 16'hFFFC;
rommem[3018] <= 16'h1784;
rommem[3019] <= 16'h4DF9;
rommem[3020] <= 16'hFFDC;
rommem[3021] <= 16'h0E00;
rommem[3022] <= 16'h3D7C;
rommem[3023] <= 16'h0001;
rommem[3024] <= 16'h0004;
rommem[3025] <= 16'h3D7C;
rommem[3026] <= 16'h0076;
rommem[3027] <= 16'h0006;
rommem[3028] <= 16'h3D7C;
rommem[3029] <= 16'h0090;
rommem[3030] <= 16'h0008;
rommem[3031] <= 16'h6100;
rommem[3032] <= 16'hFE9A;
rommem[3033] <= 16'h6100;
rommem[3034] <= 16'hFEDC;
rommem[3035] <= 16'h3D7C;
rommem[3036] <= 16'h0040;
rommem[3037] <= 16'h0006;
rommem[3038] <= 16'h3D7C;
rommem[3039] <= 16'h0010;
rommem[3040] <= 16'h0008;
rommem[3041] <= 16'h6100;
rommem[3042] <= 16'hFE86;
rommem[3043] <= 16'h6100;
rommem[3044] <= 16'hFEC8;
rommem[3045] <= 16'h3D40;
rommem[3046] <= 16'h0006;
rommem[3047] <= 16'h3D7C;
rommem[3048] <= 16'h0010;
rommem[3049] <= 16'h0008;
rommem[3050] <= 16'h6100;
rommem[3051] <= 16'hFE74;
rommem[3052] <= 16'h6100;
rommem[3053] <= 16'hFEB6;
rommem[3054] <= 16'h3D58;
rommem[3055] <= 16'h0006;
rommem[3056] <= 16'h3D7C;
rommem[3057] <= 16'h0010;
rommem[3058] <= 16'h0008;
rommem[3059] <= 16'h6100;
rommem[3060] <= 16'hFE62;
rommem[3061] <= 16'h6100;
rommem[3062] <= 16'hFEA4;
rommem[3063] <= 16'h3D58;
rommem[3064] <= 16'h0006;
rommem[3065] <= 16'h3D7C;
rommem[3066] <= 16'h0010;
rommem[3067] <= 16'h0008;
rommem[3068] <= 16'h6100;
rommem[3069] <= 16'hFE50;
rommem[3070] <= 16'h6100;
rommem[3071] <= 16'hFE92;
rommem[3072] <= 16'h3D58;
rommem[3073] <= 16'h0006;
rommem[3074] <= 16'h3D7C;
rommem[3075] <= 16'h0010;
rommem[3076] <= 16'h0008;
rommem[3077] <= 16'h6100;
rommem[3078] <= 16'hFE3E;
rommem[3079] <= 16'h6100;
rommem[3080] <= 16'hFE80;
rommem[3081] <= 16'h3D58;
rommem[3082] <= 16'h0006;
rommem[3083] <= 16'h3D7C;
rommem[3084] <= 16'h0010;
rommem[3085] <= 16'h0008;
rommem[3086] <= 16'h6100;
rommem[3087] <= 16'hFE2C;
rommem[3088] <= 16'h6100;
rommem[3089] <= 16'hFE6E;
rommem[3090] <= 16'h3D58;
rommem[3091] <= 16'h0006;
rommem[3092] <= 16'h3D7C;
rommem[3093] <= 16'h0010;
rommem[3094] <= 16'h0008;
rommem[3095] <= 16'h6100;
rommem[3096] <= 16'hFE1A;
rommem[3097] <= 16'h6100;
rommem[3098] <= 16'hFE5C;
rommem[3099] <= 16'h3D58;
rommem[3100] <= 16'h0006;
rommem[3101] <= 16'h3D7C;
rommem[3102] <= 16'h0050;
rommem[3103] <= 16'h0008;
rommem[3104] <= 16'h6100;
rommem[3105] <= 16'hFE08;
rommem[3106] <= 16'h6100;
rommem[3107] <= 16'hFE4A;
rommem[3108] <= 16'h4E75;
rommem[3109] <= 16'h7021;
rommem[3110] <= 16'h7200;
rommem[3111] <= 16'h6100;
rommem[3112] <= 16'hFEDA;
rommem[3113] <= 16'h7020;
rommem[3114] <= 16'h6100;
rommem[3115] <= 16'hFED4;
rommem[3116] <= 16'h7023;
rommem[3117] <= 16'h323C;
rommem[3118] <= 16'h00E7;
rommem[3119] <= 16'h6100;
rommem[3120] <= 16'hFECA;
rommem[3121] <= 16'h7024;
rommem[3122] <= 16'h323C;
rommem[3123] <= 16'h00E7;
rommem[3124] <= 16'h6100;
rommem[3125] <= 16'hFEC0;
rommem[3126] <= 16'h4E75;
rommem[3127] <= 16'h2C7C;
rommem[3128] <= 16'hFFDC;
rommem[3129] <= 16'h0E10;
rommem[3130] <= 16'h4BF9;
rommem[3131] <= 16'h0001;
rommem[3132] <= 16'h0600;
rommem[3133] <= 16'h3D7C;
rommem[3134] <= 16'h0080;
rommem[3135] <= 16'h0004;
rommem[3136] <= 16'h303C;
rommem[3137] <= 16'h00DE;
rommem[3138] <= 16'h323C;
rommem[3139] <= 16'h0090;
rommem[3140] <= 16'h6100;
rommem[3141] <= 16'hFDD0;
rommem[3142] <= 16'h4A00;
rommem[3143] <= 16'h6B72;
rommem[3144] <= 16'h303C;
rommem[3145] <= 16'h0000;
rommem[3146] <= 16'h323C;
rommem[3147] <= 16'h0010;
rommem[3148] <= 16'h6100;
rommem[3149] <= 16'hFDC0;
rommem[3150] <= 16'h4A00;
rommem[3151] <= 16'h6B62;
rommem[3152] <= 16'h303C;
rommem[3153] <= 16'h00DF;
rommem[3154] <= 16'h323C;
rommem[3155] <= 16'h0090;
rommem[3156] <= 16'h6100;
rommem[3157] <= 16'hFDB0;
rommem[3158] <= 16'h4A00;
rommem[3159] <= 16'h6B52;
rommem[3160] <= 16'h343C;
rommem[3161] <= 16'h0020;
rommem[3162] <= 16'h3D7C;
rommem[3163] <= 16'h0020;
rommem[3164] <= 16'h0008;
rommem[3165] <= 16'h6100;
rommem[3166] <= 16'hFD8E;
rommem[3167] <= 16'h6100;
rommem[3168] <= 16'hFDD0;
rommem[3169] <= 16'h302E;
rommem[3170] <= 16'h000A;
rommem[3171] <= 16'h4A00;
rommem[3172] <= 16'h6B38;
rommem[3173] <= 16'h302E;
rommem[3174] <= 16'h0006;
rommem[3175] <= 16'h1B80;
rommem[3176] <= 16'h2000;
rommem[3177] <= 16'h5242;
rommem[3178] <= 16'hB47C;
rommem[3179] <= 16'h005F;
rommem[3180] <= 16'h66DA;
rommem[3181] <= 16'h3D7C;
rommem[3182] <= 16'h0068;
rommem[3183] <= 16'h0008;
rommem[3184] <= 16'h6100;
rommem[3185] <= 16'hFD68;
rommem[3186] <= 16'h6100;
rommem[3187] <= 16'hFDAA;
rommem[3188] <= 16'h302E;
rommem[3189] <= 16'h000A;
rommem[3190] <= 16'h4A00;
rommem[3191] <= 16'h6B12;
rommem[3192] <= 16'h302E;
rommem[3193] <= 16'h0006;
rommem[3194] <= 16'h1B80;
rommem[3195] <= 16'h2000;
rommem[3196] <= 16'h3D7C;
rommem[3197] <= 16'h0000;
rommem[3198] <= 16'h0004;
rommem[3199] <= 16'h7000;
rommem[3200] <= 16'h4E75;
rommem[3201] <= 16'h3D7C;
rommem[3202] <= 16'h0000;
rommem[3203] <= 16'h0004;
rommem[3204] <= 16'h4E75;
rommem[3205] <= 16'h2C7C;
rommem[3206] <= 16'hFFDC;
rommem[3207] <= 16'h0E10;
rommem[3208] <= 16'h4BF9;
rommem[3209] <= 16'h0001;
rommem[3210] <= 16'h0600;
rommem[3211] <= 16'h3D7C;
rommem[3212] <= 16'h0080;
rommem[3213] <= 16'h0004;
rommem[3214] <= 16'h303C;
rommem[3215] <= 16'h00DE;
rommem[3216] <= 16'h323C;
rommem[3217] <= 16'h0090;
rommem[3218] <= 16'h6100;
rommem[3219] <= 16'hFD34;
rommem[3220] <= 16'h4A00;
rommem[3221] <= 16'h6B46;
rommem[3222] <= 16'h303C;
rommem[3223] <= 16'h0000;
rommem[3224] <= 16'h323C;
rommem[3225] <= 16'h0010;
rommem[3226] <= 16'h6100;
rommem[3227] <= 16'hFD24;
rommem[3228] <= 16'h4A00;
rommem[3229] <= 16'h6B36;
rommem[3230] <= 16'h343C;
rommem[3231] <= 16'h0020;
rommem[3232] <= 16'h1035;
rommem[3233] <= 16'h2000;
rommem[3234] <= 16'h323C;
rommem[3235] <= 16'h0010;
rommem[3236] <= 16'h6100;
rommem[3237] <= 16'hFD10;
rommem[3238] <= 16'h4A00;
rommem[3239] <= 16'h6B22;
rommem[3240] <= 16'h5242;
rommem[3241] <= 16'hB47C;
rommem[3242] <= 16'h005F;
rommem[3243] <= 16'h66E8;
rommem[3244] <= 16'h1035;
rommem[3245] <= 16'h2000;
rommem[3246] <= 16'h323C;
rommem[3247] <= 16'h0050;
rommem[3248] <= 16'h6100;
rommem[3249] <= 16'hFCF8;
rommem[3250] <= 16'h4A00;
rommem[3251] <= 16'h6B0A;
rommem[3252] <= 16'h3D7C;
rommem[3253] <= 16'h0000;
rommem[3254] <= 16'h0004;
rommem[3255] <= 16'h7000;
rommem[3256] <= 16'h4E75;
rommem[3257] <= 16'h3D7C;
rommem[3258] <= 16'h0000;
rommem[3259] <= 16'h0004;
rommem[3260] <= 16'h4E75;
rommem[3261] <= 16'h5254;
rommem[3262] <= 16'h4320;
rommem[3263] <= 16'h7265;
rommem[3264] <= 16'h6164;
rommem[3265] <= 16'h2F77;
rommem[3266] <= 16'h7269;
rommem[3267] <= 16'h7465;
rommem[3268] <= 16'h2066;
rommem[3269] <= 16'h6169;
rommem[3270] <= 16'h6C65;
rommem[3271] <= 16'h642E;
rommem[3272] <= 16'h0D0A;
rommem[3273] <= 16'h00FF;
rommem[3274] <= 16'h48E7;
rommem[3275] <= 16'h8004;
rommem[3276] <= 16'h4BF9;
rommem[3277] <= 16'hFFE0;
rommem[3278] <= 16'h0000;
rommem[3279] <= 16'h2B7C;
rommem[3280] <= 16'h0000;
rommem[3281] <= 16'h0004;
rommem[3282] <= 16'h0700;
rommem[3283] <= 16'h3B7C;
rommem[3284] <= 16'h00F3;
rommem[3285] <= 16'h0708;
rommem[3286] <= 16'h202D;
rommem[3287] <= 16'h0704;
rommem[3288] <= 16'h0800;
rommem[3289] <= 16'h0000;
rommem[3290] <= 16'h66F0;
rommem[3291] <= 16'h4CDF;
rommem[3292] <= 16'h2001;
rommem[3293] <= 16'h4E75;
rommem[3294] <= 16'h6100;
rommem[3295] <= 16'hFFD6;
rommem[3296] <= 16'h4BF9;
rommem[3297] <= 16'hFFE0;
rommem[3298] <= 16'h0000;
rommem[3299] <= 16'h2B7C;
rommem[3300] <= 16'h0000;
rommem[3301] <= 16'h0014;
rommem[3302] <= 16'h0700;
rommem[3303] <= 16'h2B7C;
rommem[3304] <= 16'h0000;
rommem[3305] <= 16'h0190;
rommem[3306] <= 16'h0704;
rommem[3307] <= 16'h3B7C;
rommem[3308] <= 16'h00F7;
rommem[3309] <= 16'h0708;
rommem[3310] <= 16'h2B7C;
rommem[3311] <= 16'h0000;
rommem[3312] <= 16'h0018;
rommem[3313] <= 16'h0700;
rommem[3314] <= 16'h2B7C;
rommem[3315] <= 16'h0000;
rommem[3316] <= 16'h012C;
rommem[3317] <= 16'h0704;
rommem[3318] <= 16'h3B7C;
rommem[3319] <= 16'h00F7;
rommem[3320] <= 16'h0708;
rommem[3321] <= 16'h4E75;
rommem[3322] <= 16'h6100;
rommem[3323] <= 16'hFF9E;
rommem[3324] <= 16'h4BF9;
rommem[3325] <= 16'hFFE0;
rommem[3326] <= 16'h0000;
rommem[3327] <= 16'h2B7C;
rommem[3328] <= 16'h0000;
rommem[3329] <= 16'h0000;
rommem[3330] <= 16'h0700;
rommem[3331] <= 16'h23FC;
rommem[3332] <= 16'h0000;
rommem[3333] <= 16'h0000;
rommem[3334] <= 16'h0001;
rommem[3335] <= 16'h042C;
rommem[3336] <= 16'h2B7C;
rommem[3337] <= 16'h0000;
rommem[3338] <= 16'h0000;
rommem[3339] <= 16'h0704;
rommem[3340] <= 16'h3B7C;
rommem[3341] <= 16'h00F7;
rommem[3342] <= 16'h0708;
rommem[3343] <= 16'h2B7C;
rommem[3344] <= 16'h0000;
rommem[3345] <= 16'h0010;
rommem[3346] <= 16'h0700;
rommem[3347] <= 16'h3B7C;
rommem[3348] <= 16'h00F7;
rommem[3349] <= 16'h0708;
rommem[3350] <= 16'h4E75;
rommem[3351] <= 16'h4BF9;
rommem[3352] <= 16'hFFE0;
rommem[3353] <= 16'h0000;
rommem[3354] <= 16'h02B9;
rommem[3355] <= 16'hFFFF;
rommem[3356] <= 16'hFFFD;
rommem[3357] <= 16'h0001;
rommem[3358] <= 16'h042C;
rommem[3359] <= 16'h00B9;
rommem[3360] <= 16'h0000;
rommem[3361] <= 16'h0001;
rommem[3362] <= 16'h0001;
rommem[3363] <= 16'h042C;
rommem[3364] <= 16'h6100;
rommem[3365] <= 16'hFF4A;
rommem[3366] <= 16'h2B7C;
rommem[3367] <= 16'h0000;
rommem[3368] <= 16'h0000;
rommem[3369] <= 16'h0700;
rommem[3370] <= 16'h2B79;
rommem[3371] <= 16'h0001;
rommem[3372] <= 16'h042C;
rommem[3373] <= 16'h0704;
rommem[3374] <= 16'h3B7C;
rommem[3375] <= 16'h00F7;
rommem[3376] <= 16'h0708;
rommem[3377] <= 16'h4E75;
rommem[3378] <= 16'h6100;
rommem[3379] <= 16'hFF2E;
rommem[3380] <= 16'h4BF9;
rommem[3381] <= 16'hFFE0;
rommem[3382] <= 16'h0000;
rommem[3383] <= 16'h2B7C;
rommem[3384] <= 16'h0000;
rommem[3385] <= 16'h0084;
rommem[3386] <= 16'h0700;
rommem[3387] <= 16'h2B40;
rommem[3388] <= 16'h0704;
rommem[3389] <= 16'h3B7C;
rommem[3390] <= 16'h00F7;
rommem[3391] <= 16'h0708;
rommem[3392] <= 16'h4E75;
rommem[3393] <= 16'h6100;
rommem[3394] <= 16'hFF10;
rommem[3395] <= 16'h4BF9;
rommem[3396] <= 16'hFFE0;
rommem[3397] <= 16'h0000;
rommem[3398] <= 16'h2B7C;
rommem[3399] <= 16'h0000;
rommem[3400] <= 16'h0038;
rommem[3401] <= 16'h0700;
rommem[3402] <= 16'h2B40;
rommem[3403] <= 16'h0704;
rommem[3404] <= 16'h3B7C;
rommem[3405] <= 16'h00F7;
rommem[3406] <= 16'h0708;
rommem[3407] <= 16'h2B7C;
rommem[3408] <= 16'h0000;
rommem[3409] <= 16'h003C;
rommem[3410] <= 16'h0700;
rommem[3411] <= 16'h2B41;
rommem[3412] <= 16'h0704;
rommem[3413] <= 16'h3B7C;
rommem[3414] <= 16'h00F7;
rommem[3415] <= 16'h0708;
rommem[3416] <= 16'h2B7C;
rommem[3417] <= 16'h0000;
rommem[3418] <= 16'h0040;
rommem[3419] <= 16'h0700;
rommem[3420] <= 16'h2B7C;
rommem[3421] <= 16'h0000;
rommem[3422] <= 16'h0000;
rommem[3423] <= 16'h0704;
rommem[3424] <= 16'h3B7C;
rommem[3425] <= 16'h00F7;
rommem[3426] <= 16'h0708;
rommem[3427] <= 16'h2C39;
rommem[3428] <= 16'h0001;
rommem[3429] <= 16'h042C;
rommem[3430] <= 16'h0086;
rommem[3431] <= 16'h0000;
rommem[3432] <= 16'h0000;
rommem[3433] <= 16'h2A86;
rommem[3434] <= 16'h2B46;
rommem[3435] <= 16'h0704;
rommem[3436] <= 16'h3B7C;
rommem[3437] <= 16'h00F7;
rommem[3438] <= 16'h0708;
rommem[3439] <= 16'h2B7C;
rommem[3440] <= 16'h0000;
rommem[3441] <= 16'h0038;
rommem[3442] <= 16'h0700;
rommem[3443] <= 16'h2B42;
rommem[3444] <= 16'h0704;
rommem[3445] <= 16'h3B7C;
rommem[3446] <= 16'h00F7;
rommem[3447] <= 16'h0708;
rommem[3448] <= 16'h2B7C;
rommem[3449] <= 16'h0000;
rommem[3450] <= 16'h003C;
rommem[3451] <= 16'h0700;
rommem[3452] <= 16'h2B43;
rommem[3453] <= 16'h0704;
rommem[3454] <= 16'h3B7C;
rommem[3455] <= 16'h00F7;
rommem[3456] <= 16'h0708;
rommem[3457] <= 16'h2B7C;
rommem[3458] <= 16'h0000;
rommem[3459] <= 16'h0040;
rommem[3460] <= 16'h0700;
rommem[3461] <= 16'h2B7C;
rommem[3462] <= 16'h0000;
rommem[3463] <= 16'h0000;
rommem[3464] <= 16'h0704;
rommem[3465] <= 16'h3B7C;
rommem[3466] <= 16'h00F7;
rommem[3467] <= 16'h0708;
rommem[3468] <= 16'h2C39;
rommem[3469] <= 16'h0001;
rommem[3470] <= 16'h042C;
rommem[3471] <= 16'h0086;
rommem[3472] <= 16'h0001;
rommem[3473] <= 16'h0000;
rommem[3474] <= 16'h2A86;
rommem[3475] <= 16'h2B46;
rommem[3476] <= 16'h0704;
rommem[3477] <= 16'h3B7C;
rommem[3478] <= 16'h00F7;
rommem[3479] <= 16'h0708;
rommem[3480] <= 16'h2C39;
rommem[3481] <= 16'h0001;
rommem[3482] <= 16'h042C;
rommem[3483] <= 16'h0086;
rommem[3484] <= 16'h0000;
rommem[3485] <= 16'h0200;
rommem[3486] <= 16'h2A86;
rommem[3487] <= 16'h2B46;
rommem[3488] <= 16'h0704;
rommem[3489] <= 16'h3B7C;
rommem[3490] <= 16'h00F7;
rommem[3491] <= 16'h0708;
rommem[3492] <= 16'h4E75;
rommem[3493] <= 16'h6100;
rommem[3494] <= 16'hFEA8;
rommem[3495] <= 16'h6100;
rommem[3496] <= 16'hFE6C;
rommem[3497] <= 16'h4DF9;
rommem[3498] <= 16'hFFDC;
rommem[3499] <= 16'h0000;
rommem[3500] <= 16'h202E;
rommem[3501] <= 16'h0C00;
rommem[3502] <= 16'h3200;
rommem[3503] <= 16'h4840;
rommem[3504] <= 16'h0240;
rommem[3505] <= 16'h00FF;
rommem[3506] <= 16'h0241;
rommem[3507] <= 16'h00FF;
rommem[3508] <= 16'h426E;
rommem[3509] <= 16'h0C04;
rommem[3510] <= 16'h242E;
rommem[3511] <= 16'h0C00;
rommem[3512] <= 16'h3602;
rommem[3513] <= 16'h4842;
rommem[3514] <= 16'h0242;
rommem[3515] <= 16'h00FF;
rommem[3516] <= 16'h0243;
rommem[3517] <= 16'h00FF;
rommem[3518] <= 16'h426E;
rommem[3519] <= 16'h0C04;
rommem[3520] <= 16'h282E;
rommem[3521] <= 16'h0C00;
rommem[3522] <= 16'h0244;
rommem[3523] <= 16'h7FFF;
rommem[3524] <= 16'h426E;
rommem[3525] <= 16'h0C04;
rommem[3526] <= 16'h2C00;
rommem[3527] <= 16'h2004;
rommem[3528] <= 16'h6100;
rommem[3529] <= 16'hFED2;
rommem[3530] <= 16'h2006;
rommem[3531] <= 16'h6100;
rommem[3532] <= 16'hFEEA;
rommem[3533] <= 16'h60B6;
rommem[3534] <= 16'h4E34;
rommem[3535] <= 16'h5620;
rommem[3536] <= 16'h3638;
rommem[3537] <= 16'h6B20;
rommem[3538] <= 16'h5379;
rommem[3539] <= 16'h7374;
rommem[3540] <= 16'h656D;
rommem[3541] <= 16'h2053;
rommem[3542] <= 16'h7461;
rommem[3543] <= 16'h7274;
rommem[3544] <= 16'h696E;
rommem[3545] <= 16'h6700;
rommem[3546] <= 16'h33FC;
rommem[3547] <= 16'h1010;
rommem[3548] <= 16'hFFDC;
rommem[3549] <= 16'h0600;
rommem[3550] <= 16'h223C;
rommem[3551] <= 16'h0002;
rommem[3552] <= 16'h0000;
rommem[3553] <= 16'h207C;
rommem[3554] <= 16'h1FF4;
rommem[3555] <= 16'h0000;
rommem[3556] <= 16'h7007;
rommem[3557] <= 16'h20C0;
rommem[3558] <= 16'h0680;
rommem[3559] <= 16'h0000;
rommem[3560] <= 16'h1000;
rommem[3561] <= 16'h5381;
rommem[3562] <= 16'h66F4;
rommem[3563] <= 16'h33FC;
rommem[3564] <= 16'h1111;
rommem[3565] <= 16'hFFDC;
rommem[3566] <= 16'h0600;
rommem[3567] <= 16'h323C;
rommem[3568] <= 16'h0400;
rommem[3569] <= 16'h207C;
rommem[3570] <= 16'h1FFF;
rommem[3571] <= 16'hE000;
rommem[3572] <= 16'h203C;
rommem[3573] <= 16'h1FFF;
rommem[3574] <= 16'hD006;
rommem[3575] <= 16'h20C0;
rommem[3576] <= 16'h51C9;
rommem[3577] <= 16'hFFFC;
rommem[3578] <= 16'h33FC;
rommem[3579] <= 16'h1212;
rommem[3580] <= 16'hFFDC;
rommem[3581] <= 16'h0600;
rommem[3582] <= 16'h747F;
rommem[3583] <= 16'h207C;
rommem[3584] <= 16'h1FFF;
rommem[3585] <= 16'hF000;
rommem[3586] <= 16'h223C;
rommem[3587] <= 16'h1FFF;
rommem[3588] <= 16'hE000;
rommem[3589] <= 16'h203C;
rommem[3590] <= 16'h1FF4;
rommem[3591] <= 16'h0007;
rommem[3592] <= 16'h2141;
rommem[3593] <= 16'h0200;
rommem[3594] <= 16'h2141;
rommem[3595] <= 16'h0400;
rommem[3596] <= 16'h2141;
rommem[3597] <= 16'h0600;
rommem[3598] <= 16'h2141;
rommem[3599] <= 16'h0800;
rommem[3600] <= 16'h2141;
rommem[3601] <= 16'h0A00;
rommem[3602] <= 16'h2141;
rommem[3603] <= 16'h0C00;
rommem[3604] <= 16'h2141;
rommem[3605] <= 16'h0E00;
rommem[3606] <= 16'h20C0;
rommem[3607] <= 16'h0680;
rommem[3608] <= 16'h0000;
rommem[3609] <= 16'h1000;
rommem[3610] <= 16'h51CA;
rommem[3611] <= 16'hFFDA;
rommem[3612] <= 16'h33FC;
rommem[3613] <= 16'h1919;
rommem[3614] <= 16'hFFDC;
rommem[3615] <= 16'h0600;
rommem[3616] <= 16'h33FC;
rommem[3617] <= 16'h0000;
rommem[3618] <= 16'hFFFF;
rommem[3619] <= 16'hFFF6;
rommem[3620] <= 16'h23F9;
rommem[3621] <= 16'h1FFF;
rommem[3622] <= 16'hF000;
rommem[3623] <= 16'hFFFF;
rommem[3624] <= 16'hFFF0;
rommem[3625] <= 16'h4E75;
rommem[3626] <= 16'h0000;
rommem[3627] <= 16'h0000;
rommem[3628] <= 16'h0000;
rommem[3629] <= 16'h0000;
rommem[3630] <= 16'h0000;
rommem[3631] <= 16'h0000;
rommem[3632] <= 16'h0000;
rommem[3633] <= 16'h0000;
rommem[3634] <= 16'h0000;
rommem[3635] <= 16'h0000;
rommem[3636] <= 16'h0000;
rommem[3637] <= 16'h0000;
rommem[3638] <= 16'h0000;
rommem[3639] <= 16'h0000;
rommem[3640] <= 16'h0000;
rommem[3641] <= 16'h0000;
rommem[3642] <= 16'h0000;
rommem[3643] <= 16'h0000;
rommem[3644] <= 16'h0000;
rommem[3645] <= 16'h0000;
rommem[3646] <= 16'h0000;
rommem[3647] <= 16'h0000;
rommem[3648] <= 16'h0000;
rommem[3649] <= 16'h0000;
rommem[3650] <= 16'h0000;
rommem[3651] <= 16'h0000;
rommem[3652] <= 16'h0000;
rommem[3653] <= 16'h0000;
rommem[3654] <= 16'h0000;
rommem[3655] <= 16'h0000;
rommem[3656] <= 16'h0000;
rommem[3657] <= 16'h0000;
rommem[3658] <= 16'h0000;
rommem[3659] <= 16'h0000;
rommem[3660] <= 16'h0000;
rommem[3661] <= 16'h0000;
rommem[3662] <= 16'h0000;
rommem[3663] <= 16'h0000;
rommem[3664] <= 16'h0000;
rommem[3665] <= 16'h0000;
rommem[3666] <= 16'h0000;
rommem[3667] <= 16'h0000;
rommem[3668] <= 16'h0000;
rommem[3669] <= 16'h0000;
rommem[3670] <= 16'h0000;
rommem[3671] <= 16'h0000;
rommem[3672] <= 16'h0000;
rommem[3673] <= 16'h0000;
rommem[3674] <= 16'h0000;
rommem[3675] <= 16'h0000;
rommem[3676] <= 16'h0000;
rommem[3677] <= 16'h0000;
rommem[3678] <= 16'h0000;
rommem[3679] <= 16'h0000;
rommem[3680] <= 16'h0000;
rommem[3681] <= 16'h0000;
rommem[3682] <= 16'h0000;
rommem[3683] <= 16'h0000;
rommem[3684] <= 16'h0000;
rommem[3685] <= 16'h0000;
rommem[3686] <= 16'h0000;
rommem[3687] <= 16'h0000;
rommem[3688] <= 16'h0000;
rommem[3689] <= 16'h0000;
rommem[3690] <= 16'h0000;
rommem[3691] <= 16'h0000;
rommem[3692] <= 16'h0000;
rommem[3693] <= 16'h0000;
rommem[3694] <= 16'h0000;
rommem[3695] <= 16'h0000;
rommem[3696] <= 16'h0000;
rommem[3697] <= 16'h0000;
rommem[3698] <= 16'h0000;
rommem[3699] <= 16'h0000;
rommem[3700] <= 16'h0000;
rommem[3701] <= 16'h0000;
rommem[3702] <= 16'h0000;
rommem[3703] <= 16'h0000;
rommem[3704] <= 16'h0000;
rommem[3705] <= 16'h0000;
rommem[3706] <= 16'h0000;
rommem[3707] <= 16'h0000;
rommem[3708] <= 16'h0000;
rommem[3709] <= 16'h0000;
rommem[3710] <= 16'h0000;
rommem[3711] <= 16'h0000;
rommem[3712] <= 16'h0000;
rommem[3713] <= 16'h0000;
rommem[3714] <= 16'h0000;
rommem[3715] <= 16'h0000;
rommem[3716] <= 16'h0000;
rommem[3717] <= 16'h0000;
rommem[3718] <= 16'h0000;
rommem[3719] <= 16'h0000;
rommem[3720] <= 16'h0000;
rommem[3721] <= 16'h0000;
rommem[3722] <= 16'h0000;
rommem[3723] <= 16'h0000;
rommem[3724] <= 16'h0000;
rommem[3725] <= 16'h0000;
rommem[3726] <= 16'h0000;
rommem[3727] <= 16'h0000;
rommem[3728] <= 16'h0000;
rommem[3729] <= 16'h0000;
rommem[3730] <= 16'h0000;
rommem[3731] <= 16'h0000;
rommem[3732] <= 16'h0000;
rommem[3733] <= 16'h0000;
rommem[3734] <= 16'h0000;
rommem[3735] <= 16'h0000;
rommem[3736] <= 16'h0000;
rommem[3737] <= 16'h0000;
rommem[3738] <= 16'h0000;
rommem[3739] <= 16'h0000;
rommem[3740] <= 16'h0000;
rommem[3741] <= 16'h0000;
rommem[3742] <= 16'h0000;
rommem[3743] <= 16'h0000;
rommem[3744] <= 16'h0000;
rommem[3745] <= 16'h0000;
rommem[3746] <= 16'h0000;
rommem[3747] <= 16'h0000;
rommem[3748] <= 16'h0000;
rommem[3749] <= 16'h0000;
rommem[3750] <= 16'h0000;
rommem[3751] <= 16'h0000;
rommem[3752] <= 16'h0000;
rommem[3753] <= 16'h0000;
rommem[3754] <= 16'h0000;
rommem[3755] <= 16'h0000;
rommem[3756] <= 16'h0000;
rommem[3757] <= 16'h0000;
rommem[3758] <= 16'h1818;
rommem[3759] <= 16'h1818;
rommem[3760] <= 16'h1800;
rommem[3761] <= 16'h1800;
rommem[3762] <= 16'h6C6C;
rommem[3763] <= 16'h0000;
rommem[3764] <= 16'h0000;
rommem[3765] <= 16'h0000;
rommem[3766] <= 16'h6C6C;
rommem[3767] <= 16'hFE6C;
rommem[3768] <= 16'hFE6C;
rommem[3769] <= 16'h6C00;
rommem[3770] <= 16'h183E;
rommem[3771] <= 16'h603C;
rommem[3772] <= 16'h067C;
rommem[3773] <= 16'h1800;
rommem[3774] <= 16'h0066;
rommem[3775] <= 16'hACD8;
rommem[3776] <= 16'h366A;
rommem[3777] <= 16'hCC00;
rommem[3778] <= 16'h386C;
rommem[3779] <= 16'h6876;
rommem[3780] <= 16'hDCCE;
rommem[3781] <= 16'h7B00;
rommem[3782] <= 16'h1818;
rommem[3783] <= 16'h3000;
rommem[3784] <= 16'h0000;
rommem[3785] <= 16'h0000;
rommem[3786] <= 16'h0C18;
rommem[3787] <= 16'h3030;
rommem[3788] <= 16'h3018;
rommem[3789] <= 16'h0C00;
rommem[3790] <= 16'h3018;
rommem[3791] <= 16'h0C0C;
rommem[3792] <= 16'h0C18;
rommem[3793] <= 16'h3000;
rommem[3794] <= 16'h0066;
rommem[3795] <= 16'h3CFF;
rommem[3796] <= 16'h3C66;
rommem[3797] <= 16'h0000;
rommem[3798] <= 16'h0018;
rommem[3799] <= 16'h187E;
rommem[3800] <= 16'h1818;
rommem[3801] <= 16'h0000;
rommem[3802] <= 16'h0000;
rommem[3803] <= 16'h0000;
rommem[3804] <= 16'h0018;
rommem[3805] <= 16'h1830;
rommem[3806] <= 16'h0000;
rommem[3807] <= 16'h007E;
rommem[3808] <= 16'h0000;
rommem[3809] <= 16'h0000;
rommem[3810] <= 16'h0000;
rommem[3811] <= 16'h0000;
rommem[3812] <= 16'h0018;
rommem[3813] <= 16'h1800;
rommem[3814] <= 16'h0306;
rommem[3815] <= 16'h0C18;
rommem[3816] <= 16'h3060;
rommem[3817] <= 16'hC000;
rommem[3818] <= 16'h3C66;
rommem[3819] <= 16'h6E7E;
rommem[3820] <= 16'h7666;
rommem[3821] <= 16'h3C00;
rommem[3822] <= 16'h1838;
rommem[3823] <= 16'h7818;
rommem[3824] <= 16'h1818;
rommem[3825] <= 16'h1800;
rommem[3826] <= 16'h3C66;
rommem[3827] <= 16'h060C;
rommem[3828] <= 16'h1830;
rommem[3829] <= 16'h7E00;
rommem[3830] <= 16'h3C66;
rommem[3831] <= 16'h061C;
rommem[3832] <= 16'h0666;
rommem[3833] <= 16'h3C00;
rommem[3834] <= 16'h1C3C;
rommem[3835] <= 16'h6CCC;
rommem[3836] <= 16'hFE0C;
rommem[3837] <= 16'h0C00;
rommem[3838] <= 16'h7E60;
rommem[3839] <= 16'h7C06;
rommem[3840] <= 16'h0666;
rommem[3841] <= 16'h3C00;
rommem[3842] <= 16'h1C30;
rommem[3843] <= 16'h607C;
rommem[3844] <= 16'h6666;
rommem[3845] <= 16'h3C00;
rommem[3846] <= 16'h7E06;
rommem[3847] <= 16'h060C;
rommem[3848] <= 16'h1818;
rommem[3849] <= 16'h1800;
rommem[3850] <= 16'h3C66;
rommem[3851] <= 16'h663C;
rommem[3852] <= 16'h6666;
rommem[3853] <= 16'h3C00;
rommem[3854] <= 16'h3C66;
rommem[3855] <= 16'h663E;
rommem[3856] <= 16'h060C;
rommem[3857] <= 16'h3800;
rommem[3858] <= 16'h0018;
rommem[3859] <= 16'h1800;
rommem[3860] <= 16'h0018;
rommem[3861] <= 16'h1800;
rommem[3862] <= 16'h0018;
rommem[3863] <= 16'h1800;
rommem[3864] <= 16'h0018;
rommem[3865] <= 16'h1830;
rommem[3866] <= 16'h0006;
rommem[3867] <= 16'h1860;
rommem[3868] <= 16'h1806;
rommem[3869] <= 16'h0000;
rommem[3870] <= 16'h0000;
rommem[3871] <= 16'h7E00;
rommem[3872] <= 16'h7E00;
rommem[3873] <= 16'h0000;
rommem[3874] <= 16'h0060;
rommem[3875] <= 16'h1806;
rommem[3876] <= 16'h1860;
rommem[3877] <= 16'h0000;
rommem[3878] <= 16'h3C66;
rommem[3879] <= 16'h060C;
rommem[3880] <= 16'h1800;
rommem[3881] <= 16'h1800;
rommem[3882] <= 16'h7CC6;
rommem[3883] <= 16'hDED6;
rommem[3884] <= 16'hDEC0;
rommem[3885] <= 16'h7800;
rommem[3886] <= 16'h3C66;
rommem[3887] <= 16'h667E;
rommem[3888] <= 16'h6666;
rommem[3889] <= 16'h6600;
rommem[3890] <= 16'h7C66;
rommem[3891] <= 16'h667C;
rommem[3892] <= 16'h6666;
rommem[3893] <= 16'h7C00;
rommem[3894] <= 16'h1E30;
rommem[3895] <= 16'h6060;
rommem[3896] <= 16'h6030;
rommem[3897] <= 16'h1E00;
rommem[3898] <= 16'h786C;
rommem[3899] <= 16'h6666;
rommem[3900] <= 16'h666C;
rommem[3901] <= 16'h7800;
rommem[3902] <= 16'h7E60;
rommem[3903] <= 16'h6078;
rommem[3904] <= 16'h6060;
rommem[3905] <= 16'h7E00;
rommem[3906] <= 16'h7E60;
rommem[3907] <= 16'h6078;
rommem[3908] <= 16'h6060;
rommem[3909] <= 16'h6000;
rommem[3910] <= 16'h3C66;
rommem[3911] <= 16'h606E;
rommem[3912] <= 16'h6666;
rommem[3913] <= 16'h3E00;
rommem[3914] <= 16'h6666;
rommem[3915] <= 16'h667E;
rommem[3916] <= 16'h6666;
rommem[3917] <= 16'h6600;
rommem[3918] <= 16'h3C18;
rommem[3919] <= 16'h1818;
rommem[3920] <= 16'h1818;
rommem[3921] <= 16'h3C00;
rommem[3922] <= 16'h0606;
rommem[3923] <= 16'h0606;
rommem[3924] <= 16'h0666;
rommem[3925] <= 16'h3C00;
rommem[3926] <= 16'hC6CC;
rommem[3927] <= 16'hD8F0;
rommem[3928] <= 16'hD8CC;
rommem[3929] <= 16'hC600;
rommem[3930] <= 16'h6060;
rommem[3931] <= 16'h6060;
rommem[3932] <= 16'h6060;
rommem[3933] <= 16'h7E00;
rommem[3934] <= 16'hC6EE;
rommem[3935] <= 16'hFED6;
rommem[3936] <= 16'hC6C6;
rommem[3937] <= 16'hC600;
rommem[3938] <= 16'hC6E6;
rommem[3939] <= 16'hF6DE;
rommem[3940] <= 16'hCEC6;
rommem[3941] <= 16'hC600;
rommem[3942] <= 16'h3C66;
rommem[3943] <= 16'h6666;
rommem[3944] <= 16'h6666;
rommem[3945] <= 16'h3C00;
rommem[3946] <= 16'h7C66;
rommem[3947] <= 16'h667C;
rommem[3948] <= 16'h6060;
rommem[3949] <= 16'h6000;
rommem[3950] <= 16'h78CC;
rommem[3951] <= 16'hCCCC;
rommem[3952] <= 16'hCCDC;
rommem[3953] <= 16'h7E00;
rommem[3954] <= 16'h7C66;
rommem[3955] <= 16'h667C;
rommem[3956] <= 16'h6C66;
rommem[3957] <= 16'h6600;
rommem[3958] <= 16'h3C66;
rommem[3959] <= 16'h703C;
rommem[3960] <= 16'h0E66;
rommem[3961] <= 16'h3C00;
rommem[3962] <= 16'h7E18;
rommem[3963] <= 16'h1818;
rommem[3964] <= 16'h1818;
rommem[3965] <= 16'h1800;
rommem[3966] <= 16'h6666;
rommem[3967] <= 16'h6666;
rommem[3968] <= 16'h6666;
rommem[3969] <= 16'h3C00;
rommem[3970] <= 16'h6666;
rommem[3971] <= 16'h6666;
rommem[3972] <= 16'h3C3C;
rommem[3973] <= 16'h1800;
rommem[3974] <= 16'hC6C6;
rommem[3975] <= 16'hC6D6;
rommem[3976] <= 16'hFEEE;
rommem[3977] <= 16'hC600;
rommem[3978] <= 16'hC366;
rommem[3979] <= 16'h3C18;
rommem[3980] <= 16'h3C66;
rommem[3981] <= 16'hC300;
rommem[3982] <= 16'hC366;
rommem[3983] <= 16'h3C18;
rommem[3984] <= 16'h1818;
rommem[3985] <= 16'h1800;
rommem[3986] <= 16'hFE0C;
rommem[3987] <= 16'h1830;
rommem[3988] <= 16'h60C0;
rommem[3989] <= 16'hFE00;
rommem[3990] <= 16'h3C30;
rommem[3991] <= 16'h3030;
rommem[3992] <= 16'h3030;
rommem[3993] <= 16'h3C00;
rommem[3994] <= 16'hC060;
rommem[3995] <= 16'h3018;
rommem[3996] <= 16'h0C06;
rommem[3997] <= 16'h0300;
rommem[3998] <= 16'h3C0C;
rommem[3999] <= 16'h0C0C;
rommem[4000] <= 16'h0C0C;
rommem[4001] <= 16'h3C00;
rommem[4002] <= 16'h1038;
rommem[4003] <= 16'h6CC6;
rommem[4004] <= 16'h0000;
rommem[4005] <= 16'h0000;
rommem[4006] <= 16'h0000;
rommem[4007] <= 16'h0000;
rommem[4008] <= 16'h0000;
rommem[4009] <= 16'h00FE;
rommem[4010] <= 16'h1818;
rommem[4011] <= 16'h0C00;
rommem[4012] <= 16'h0000;
rommem[4013] <= 16'h0000;
rommem[4014] <= 16'h0000;
rommem[4015] <= 16'h3C06;
rommem[4016] <= 16'h3E66;
rommem[4017] <= 16'h3E00;
rommem[4018] <= 16'h6060;
rommem[4019] <= 16'h7C66;
rommem[4020] <= 16'h6666;
rommem[4021] <= 16'h7C00;
rommem[4022] <= 16'h0000;
rommem[4023] <= 16'h3C60;
rommem[4024] <= 16'h6060;
rommem[4025] <= 16'h3C00;
rommem[4026] <= 16'h0606;
rommem[4027] <= 16'h3E66;
rommem[4028] <= 16'h6666;
rommem[4029] <= 16'h3E00;
rommem[4030] <= 16'h0000;
rommem[4031] <= 16'h3C66;
rommem[4032] <= 16'h7E60;
rommem[4033] <= 16'h3C00;
rommem[4034] <= 16'h1C30;
rommem[4035] <= 16'h7C30;
rommem[4036] <= 16'h3030;
rommem[4037] <= 16'h3000;
rommem[4038] <= 16'h0000;
rommem[4039] <= 16'h3E66;
rommem[4040] <= 16'h663E;
rommem[4041] <= 16'h063C;
rommem[4042] <= 16'h6060;
rommem[4043] <= 16'h7C66;
rommem[4044] <= 16'h6666;
rommem[4045] <= 16'h6600;
rommem[4046] <= 16'h1800;
rommem[4047] <= 16'h1818;
rommem[4048] <= 16'h1818;
rommem[4049] <= 16'h0C00;
rommem[4050] <= 16'h0C00;
rommem[4051] <= 16'h0C0C;
rommem[4052] <= 16'h0C0C;
rommem[4053] <= 16'h0C78;
rommem[4054] <= 16'h6060;
rommem[4055] <= 16'h666C;
rommem[4056] <= 16'h786C;
rommem[4057] <= 16'h6600;
rommem[4058] <= 16'h1818;
rommem[4059] <= 16'h1818;
rommem[4060] <= 16'h1818;
rommem[4061] <= 16'h0C00;
rommem[4062] <= 16'h0000;
rommem[4063] <= 16'hECFE;
rommem[4064] <= 16'hD6C6;
rommem[4065] <= 16'hC600;
rommem[4066] <= 16'h0000;
rommem[4067] <= 16'h7C66;
rommem[4068] <= 16'h6666;
rommem[4069] <= 16'h6600;
rommem[4070] <= 16'h0000;
rommem[4071] <= 16'h3C66;
rommem[4072] <= 16'h6666;
rommem[4073] <= 16'h3C00;
rommem[4074] <= 16'h0000;
rommem[4075] <= 16'h7C66;
rommem[4076] <= 16'h667C;
rommem[4077] <= 16'h6060;
rommem[4078] <= 16'h0000;
rommem[4079] <= 16'h3E66;
rommem[4080] <= 16'h663E;
rommem[4081] <= 16'h0606;
rommem[4082] <= 16'h0000;
rommem[4083] <= 16'h7C66;
rommem[4084] <= 16'h6060;
rommem[4085] <= 16'h6000;
rommem[4086] <= 16'h0000;
rommem[4087] <= 16'h3C60;
rommem[4088] <= 16'h3C06;
rommem[4089] <= 16'h7C00;
rommem[4090] <= 16'h3030;
rommem[4091] <= 16'h7C30;
rommem[4092] <= 16'h3030;
rommem[4093] <= 16'h1C00;
rommem[4094] <= 16'h0000;
rommem[4095] <= 16'h6666;
rommem[4096] <= 16'h6666;
rommem[4097] <= 16'h3E00;
rommem[4098] <= 16'h0000;
rommem[4099] <= 16'h6666;
rommem[4100] <= 16'h663C;
rommem[4101] <= 16'h1800;
rommem[4102] <= 16'h0000;
rommem[4103] <= 16'hC6C6;
rommem[4104] <= 16'hD6FE;
rommem[4105] <= 16'h6C00;
rommem[4106] <= 16'h0000;
rommem[4107] <= 16'hC66C;
rommem[4108] <= 16'h386C;
rommem[4109] <= 16'hC600;
rommem[4110] <= 16'h0000;
rommem[4111] <= 16'h6666;
rommem[4112] <= 16'h663C;
rommem[4113] <= 16'h1830;
rommem[4114] <= 16'h0000;
rommem[4115] <= 16'h7E0C;
rommem[4116] <= 16'h1830;
rommem[4117] <= 16'h7E00;
rommem[4118] <= 16'h0E18;
rommem[4119] <= 16'h1870;
rommem[4120] <= 16'h1818;
rommem[4121] <= 16'h0E00;
rommem[4122] <= 16'h1818;
rommem[4123] <= 16'h1818;
rommem[4124] <= 16'h1818;
rommem[4125] <= 16'h1800;
rommem[4126] <= 16'h7018;
rommem[4127] <= 16'h180E;
rommem[4128] <= 16'h1818;
rommem[4129] <= 16'h7000;
rommem[4130] <= 16'h729C;
rommem[4131] <= 16'h0000;
rommem[4132] <= 16'h0000;
rommem[4133] <= 16'h0000;
rommem[4134] <= 16'hFEFE;
rommem[4135] <= 16'hFEFE;
rommem[4136] <= 16'hFEFE;
rommem[4137] <= 16'hFE00;
rommem[4138] <= 16'h0000;
rommem[4139] <= 16'h0000;
rommem[4140] <= 16'h0000;
rommem[4141] <= 16'h0000;
rommem[4142] <= 16'h0000;
rommem[4143] <= 16'h0000;
rommem[4144] <= 16'h0000;
rommem[4145] <= 16'h0000;
rommem[4146] <= 16'h0000;
rommem[4147] <= 16'h0000;
rommem[4148] <= 16'h0000;
rommem[4149] <= 16'h0000;
rommem[4150] <= 16'h0000;
rommem[4151] <= 16'h0000;
rommem[4152] <= 16'h0000;
rommem[4153] <= 16'h0000;
rommem[4154] <= 16'h0000;
rommem[4155] <= 16'h0000;
rommem[4156] <= 16'h0000;
rommem[4157] <= 16'h0000;
rommem[4158] <= 16'h0000;
rommem[4159] <= 16'h0000;
rommem[4160] <= 16'h0000;
rommem[4161] <= 16'h0000;
rommem[4162] <= 16'h0000;
rommem[4163] <= 16'h0000;
rommem[4164] <= 16'h0000;
rommem[4165] <= 16'h0000;
rommem[4166] <= 16'h0000;
rommem[4167] <= 16'h0000;
rommem[4168] <= 16'h0000;
rommem[4169] <= 16'h0000;
rommem[4170] <= 16'h0000;
rommem[4171] <= 16'h0000;
rommem[4172] <= 16'h0000;
rommem[4173] <= 16'h0000;
rommem[4174] <= 16'h0000;
rommem[4175] <= 16'h0000;
rommem[4176] <= 16'h0000;
rommem[4177] <= 16'h0000;
rommem[4178] <= 16'h0000;
rommem[4179] <= 16'h0000;
rommem[4180] <= 16'h0000;
rommem[4181] <= 16'h0000;
rommem[4182] <= 16'h0000;
rommem[4183] <= 16'h0000;
rommem[4184] <= 16'h0000;
rommem[4185] <= 16'h0000;
rommem[4186] <= 16'h0000;
rommem[4187] <= 16'h0000;
rommem[4188] <= 16'h0000;
rommem[4189] <= 16'h0000;
rommem[4190] <= 16'h0000;
rommem[4191] <= 16'h0000;
rommem[4192] <= 16'h0000;
rommem[4193] <= 16'h0000;
rommem[4194] <= 16'h0000;
rommem[4195] <= 16'h0000;
rommem[4196] <= 16'h0000;
rommem[4197] <= 16'h0000;
rommem[4198] <= 16'h0000;
rommem[4199] <= 16'h0000;
rommem[4200] <= 16'h0000;
rommem[4201] <= 16'h0000;
rommem[4202] <= 16'h0000;
rommem[4203] <= 16'h0000;
rommem[4204] <= 16'h0000;
rommem[4205] <= 16'h0000;
rommem[4206] <= 16'h0000;
rommem[4207] <= 16'h0000;
rommem[4208] <= 16'h0000;
rommem[4209] <= 16'h0000;
rommem[4210] <= 16'h0000;
rommem[4211] <= 16'h0000;
rommem[4212] <= 16'h0000;
rommem[4213] <= 16'h0000;
rommem[4214] <= 16'h0000;
rommem[4215] <= 16'h0000;
rommem[4216] <= 16'h0000;
rommem[4217] <= 16'h0000;
rommem[4218] <= 16'h0000;
rommem[4219] <= 16'h0000;
rommem[4220] <= 16'h0000;
rommem[4221] <= 16'h0000;
rommem[4222] <= 16'h0000;
rommem[4223] <= 16'h0000;
rommem[4224] <= 16'h0000;
rommem[4225] <= 16'h0000;
rommem[4226] <= 16'h0000;
rommem[4227] <= 16'h0000;
rommem[4228] <= 16'h0000;
rommem[4229] <= 16'h0000;
rommem[4230] <= 16'h0000;
rommem[4231] <= 16'h0000;
rommem[4232] <= 16'h0000;
rommem[4233] <= 16'h0000;
rommem[4234] <= 16'h0000;
rommem[4235] <= 16'h0000;
rommem[4236] <= 16'h0000;
rommem[4237] <= 16'h0000;
rommem[4238] <= 16'h0000;
rommem[4239] <= 16'h0000;
rommem[4240] <= 16'h0000;
rommem[4241] <= 16'h0000;
rommem[4242] <= 16'h0000;
rommem[4243] <= 16'h0000;
rommem[4244] <= 16'h0000;
rommem[4245] <= 16'h0000;
rommem[4246] <= 16'h0000;
rommem[4247] <= 16'h0000;
rommem[4248] <= 16'h0000;
rommem[4249] <= 16'h0000;
rommem[4250] <= 16'h0000;
rommem[4251] <= 16'h0000;
rommem[4252] <= 16'h0000;
rommem[4253] <= 16'h0000;
rommem[4254] <= 16'h0000;
rommem[4255] <= 16'h0000;
rommem[4256] <= 16'h0000;
rommem[4257] <= 16'h0000;
rommem[4258] <= 16'h0000;
rommem[4259] <= 16'h0000;
rommem[4260] <= 16'h0000;
rommem[4261] <= 16'h0000;
rommem[4262] <= 16'h0000;
rommem[4263] <= 16'h0000;
rommem[4264] <= 16'h0000;
rommem[4265] <= 16'h0000;
rommem[4266] <= 16'h0000;
rommem[4267] <= 16'h0000;
rommem[4268] <= 16'h0000;
rommem[4269] <= 16'h0000;
rommem[4270] <= 16'h0000;
rommem[4271] <= 16'h0000;
rommem[4272] <= 16'h0000;
rommem[4273] <= 16'h0000;
rommem[4274] <= 16'h0000;
rommem[4275] <= 16'h0000;
rommem[4276] <= 16'h0000;
rommem[4277] <= 16'h0000;
rommem[4278] <= 16'h0000;
rommem[4279] <= 16'h0000;
rommem[4280] <= 16'h0000;
rommem[4281] <= 16'h0000;
rommem[4282] <= 16'h0000;
rommem[4283] <= 16'h0000;
rommem[4284] <= 16'h0000;
rommem[4285] <= 16'h0000;
rommem[4286] <= 16'h0000;
rommem[4287] <= 16'h0000;
rommem[4288] <= 16'h0000;
rommem[4289] <= 16'h0000;
rommem[4290] <= 16'h0000;
rommem[4291] <= 16'h0000;
rommem[4292] <= 16'h0000;
rommem[4293] <= 16'h0000;
rommem[4294] <= 16'h0000;
rommem[4295] <= 16'h0000;
rommem[4296] <= 16'h0000;
rommem[4297] <= 16'h0000;
rommem[4298] <= 16'h0000;
rommem[4299] <= 16'h0000;
rommem[4300] <= 16'h0000;
rommem[4301] <= 16'h0000;
rommem[4302] <= 16'h0000;
rommem[4303] <= 16'h0000;
rommem[4304] <= 16'h0000;
rommem[4305] <= 16'h0000;
rommem[4306] <= 16'h0000;
rommem[4307] <= 16'h0000;
rommem[4308] <= 16'h0000;
rommem[4309] <= 16'h0000;
rommem[4310] <= 16'h0000;
rommem[4311] <= 16'h0000;
rommem[4312] <= 16'h0000;
rommem[4313] <= 16'h0000;
rommem[4314] <= 16'h0000;
rommem[4315] <= 16'h0000;
rommem[4316] <= 16'h0000;
rommem[4317] <= 16'h0000;
rommem[4318] <= 16'h0000;
rommem[4319] <= 16'h0000;
rommem[4320] <= 16'h0000;
rommem[4321] <= 16'h0000;
rommem[4322] <= 16'h0000;
rommem[4323] <= 16'h0000;
rommem[4324] <= 16'h0000;
rommem[4325] <= 16'h0000;
rommem[4326] <= 16'h0000;
rommem[4327] <= 16'h0000;
rommem[4328] <= 16'h0000;
rommem[4329] <= 16'h0000;
rommem[4330] <= 16'h0000;
rommem[4331] <= 16'h0000;
rommem[4332] <= 16'h0000;
rommem[4333] <= 16'h0000;
rommem[4334] <= 16'h0000;
rommem[4335] <= 16'h0000;
rommem[4336] <= 16'h0000;
rommem[4337] <= 16'h0000;
rommem[4338] <= 16'h0000;
rommem[4339] <= 16'h0000;
rommem[4340] <= 16'h0000;
rommem[4341] <= 16'h0000;
rommem[4342] <= 16'h0000;
rommem[4343] <= 16'h0000;
rommem[4344] <= 16'h0000;
rommem[4345] <= 16'h0000;
rommem[4346] <= 16'h0000;
rommem[4347] <= 16'h0000;
rommem[4348] <= 16'h0000;
rommem[4349] <= 16'h0000;
rommem[4350] <= 16'h0000;
rommem[4351] <= 16'h0000;
rommem[4352] <= 16'h0000;
rommem[4353] <= 16'h0000;
rommem[4354] <= 16'h0000;
rommem[4355] <= 16'h0000;
rommem[4356] <= 16'h0000;
rommem[4357] <= 16'h0000;
rommem[4358] <= 16'h0000;
rommem[4359] <= 16'h0000;
rommem[4360] <= 16'h0000;
rommem[4361] <= 16'h0000;
rommem[4362] <= 16'h0000;
rommem[4363] <= 16'h0000;
rommem[4364] <= 16'h0000;
rommem[4365] <= 16'h0000;
rommem[4366] <= 16'h0000;
rommem[4367] <= 16'h0000;
rommem[4368] <= 16'h0000;
rommem[4369] <= 16'h0000;
rommem[4370] <= 16'h0000;
rommem[4371] <= 16'h0000;
rommem[4372] <= 16'h0000;
rommem[4373] <= 16'h0000;
rommem[4374] <= 16'h0000;
rommem[4375] <= 16'h0000;
rommem[4376] <= 16'h0000;
rommem[4377] <= 16'h0000;
rommem[4378] <= 16'h0000;
rommem[4379] <= 16'h0000;
rommem[4380] <= 16'h0000;
rommem[4381] <= 16'h0000;
rommem[4382] <= 16'h0000;
rommem[4383] <= 16'h0000;
rommem[4384] <= 16'h0000;
rommem[4385] <= 16'h0000;
rommem[4386] <= 16'h0000;
rommem[4387] <= 16'h0000;
rommem[4388] <= 16'h0000;
rommem[4389] <= 16'h0000;
rommem[4390] <= 16'h0000;
rommem[4391] <= 16'h0000;
rommem[4392] <= 16'h0000;
rommem[4393] <= 16'h0000;
rommem[4394] <= 16'h0000;
rommem[4395] <= 16'h0000;
rommem[4396] <= 16'h0000;
rommem[4397] <= 16'h0000;
rommem[4398] <= 16'h0000;
rommem[4399] <= 16'h0000;
rommem[4400] <= 16'h0000;
rommem[4401] <= 16'h0000;
rommem[4402] <= 16'h0000;
rommem[4403] <= 16'h0000;
rommem[4404] <= 16'h0000;
rommem[4405] <= 16'h0000;
rommem[4406] <= 16'h0000;
rommem[4407] <= 16'h0000;
rommem[4408] <= 16'h0000;
rommem[4409] <= 16'h0000;
rommem[4410] <= 16'h0000;
rommem[4411] <= 16'h0000;
rommem[4412] <= 16'h0000;
rommem[4413] <= 16'h0000;
rommem[4414] <= 16'h0000;
rommem[4415] <= 16'h0000;
rommem[4416] <= 16'h0000;
rommem[4417] <= 16'h0000;
rommem[4418] <= 16'h0000;
rommem[4419] <= 16'h0000;
rommem[4420] <= 16'h0000;
rommem[4421] <= 16'h0000;
rommem[4422] <= 16'h0000;
rommem[4423] <= 16'h0000;
rommem[4424] <= 16'h0000;
rommem[4425] <= 16'h0000;
rommem[4426] <= 16'h0000;
rommem[4427] <= 16'h0000;
rommem[4428] <= 16'h0000;
rommem[4429] <= 16'h0000;
rommem[4430] <= 16'h0000;
rommem[4431] <= 16'h0000;
rommem[4432] <= 16'h0000;
rommem[4433] <= 16'h0000;
rommem[4434] <= 16'h0000;
rommem[4435] <= 16'h0000;
rommem[4436] <= 16'h0000;
rommem[4437] <= 16'h0000;
rommem[4438] <= 16'h0000;
rommem[4439] <= 16'h0000;
rommem[4440] <= 16'h0000;
rommem[4441] <= 16'h0000;
rommem[4442] <= 16'h0000;
rommem[4443] <= 16'h0000;
rommem[4444] <= 16'h0000;
rommem[4445] <= 16'h0000;
rommem[4446] <= 16'h0000;
rommem[4447] <= 16'h0000;
rommem[4448] <= 16'h0000;
rommem[4449] <= 16'h0000;
rommem[4450] <= 16'h0000;
rommem[4451] <= 16'h0000;
rommem[4452] <= 16'h0000;
rommem[4453] <= 16'h0000;
rommem[4454] <= 16'h0000;
rommem[4455] <= 16'h0000;
rommem[4456] <= 16'h0000;
rommem[4457] <= 16'h0000;
rommem[4458] <= 16'h0000;
rommem[4459] <= 16'h0000;
rommem[4460] <= 16'h0000;
rommem[4461] <= 16'h0000;
rommem[4462] <= 16'h0000;
rommem[4463] <= 16'h0000;
rommem[4464] <= 16'h0000;
rommem[4465] <= 16'h0000;
rommem[4466] <= 16'h0000;
rommem[4467] <= 16'h0000;
rommem[4468] <= 16'h0000;
rommem[4469] <= 16'h0000;
rommem[4470] <= 16'h0000;
rommem[4471] <= 16'h0000;
rommem[4472] <= 16'h0000;
rommem[4473] <= 16'h0000;
rommem[4474] <= 16'h0000;
rommem[4475] <= 16'h0000;
rommem[4476] <= 16'h0000;
rommem[4477] <= 16'h0000;
rommem[4478] <= 16'h0000;
rommem[4479] <= 16'h0000;
rommem[4480] <= 16'h0000;
rommem[4481] <= 16'h0000;
rommem[4482] <= 16'h0000;
rommem[4483] <= 16'h0000;
rommem[4484] <= 16'h0000;
rommem[4485] <= 16'h0000;
rommem[4486] <= 16'h0000;
rommem[4487] <= 16'h0000;
rommem[4488] <= 16'h0000;
rommem[4489] <= 16'h0000;
rommem[4490] <= 16'h0000;
rommem[4491] <= 16'h0000;
rommem[4492] <= 16'h0000;
rommem[4493] <= 16'h0000;
rommem[4494] <= 16'h0000;
rommem[4495] <= 16'h0000;
rommem[4496] <= 16'h0000;
rommem[4497] <= 16'h0000;
rommem[4498] <= 16'h0000;
rommem[4499] <= 16'h0000;
rommem[4500] <= 16'h0000;
rommem[4501] <= 16'h0000;
rommem[4502] <= 16'h0000;
rommem[4503] <= 16'h0000;
rommem[4504] <= 16'h0000;
rommem[4505] <= 16'h0000;
rommem[4506] <= 16'h0000;
rommem[4507] <= 16'h0000;
rommem[4508] <= 16'h0000;
rommem[4509] <= 16'h0000;
rommem[4510] <= 16'h0000;
rommem[4511] <= 16'h0000;
rommem[4512] <= 16'h0000;
rommem[4513] <= 16'h0000;
rommem[4514] <= 16'h0000;
rommem[4515] <= 16'h0000;
rommem[4516] <= 16'h0000;
rommem[4517] <= 16'h0000;
rommem[4518] <= 16'h0000;
rommem[4519] <= 16'h0000;
rommem[4520] <= 16'h0000;
rommem[4521] <= 16'h0000;
rommem[4522] <= 16'h0000;
rommem[4523] <= 16'h0000;
rommem[4524] <= 16'h0000;
rommem[4525] <= 16'h0000;
rommem[4526] <= 16'h0000;
rommem[4527] <= 16'h0000;
rommem[4528] <= 16'h0000;
rommem[4529] <= 16'h0000;
rommem[4530] <= 16'h0000;
rommem[4531] <= 16'h0000;
rommem[4532] <= 16'h0000;
rommem[4533] <= 16'h0000;
rommem[4534] <= 16'h0000;
rommem[4535] <= 16'h0300;
rommem[4536] <= 16'h0300;
rommem[4537] <= 16'h0300;
rommem[4538] <= 16'h0300;
rommem[4539] <= 16'h0300;
rommem[4540] <= 16'h0000;
rommem[4541] <= 16'h0300;
rommem[4542] <= 16'h0300;
rommem[4543] <= 16'h0000;
rommem[4544] <= 16'h0000;
rommem[4545] <= 16'h0000;
rommem[4546] <= 16'h0000;
rommem[4547] <= 16'h0C30;
rommem[4548] <= 16'h0C30;
rommem[4549] <= 16'h0000;
rommem[4550] <= 16'h0000;
rommem[4551] <= 16'h0000;
rommem[4552] <= 16'h0000;
rommem[4553] <= 16'h0000;
rommem[4554] <= 16'h0000;
rommem[4555] <= 16'h0000;
rommem[4556] <= 16'h0000;
rommem[4557] <= 16'h0000;
rommem[4558] <= 16'h0000;
rommem[4559] <= 16'h0C30;
rommem[4560] <= 16'h0C30;
rommem[4561] <= 16'h3FFC;
rommem[4562] <= 16'h0C30;
rommem[4563] <= 16'h0C30;
rommem[4564] <= 16'h3FFC;
rommem[4565] <= 16'h0C30;
rommem[4566] <= 16'h0C30;
rommem[4567] <= 16'h0000;
rommem[4568] <= 16'h0000;
rommem[4569] <= 16'h0000;
rommem[4570] <= 16'h0000;
rommem[4571] <= 16'h0180;
rommem[4572] <= 16'h07E0;
rommem[4573] <= 16'h0990;
rommem[4574] <= 16'h0980;
rommem[4575] <= 16'h07E0;
rommem[4576] <= 16'h0190;
rommem[4577] <= 16'h0990;
rommem[4578] <= 16'h07E0;
rommem[4579] <= 16'h0180;
rommem[4580] <= 16'h0000;
rommem[4581] <= 16'h0000;
rommem[4582] <= 16'h0000;
rommem[4583] <= 16'h0C18;
rommem[4584] <= 16'h1230;
rommem[4585] <= 16'h0C60;
rommem[4586] <= 16'h00C0;
rommem[4587] <= 16'h0180;
rommem[4588] <= 16'h0330;
rommem[4589] <= 16'h0648;
rommem[4590] <= 16'h0C30;
rommem[4591] <= 16'h0000;
rommem[4592] <= 16'h0000;
rommem[4593] <= 16'h0000;
rommem[4594] <= 16'h0000;
rommem[4595] <= 16'h0000;
rommem[4596] <= 16'h0000;
rommem[4597] <= 16'h0000;
rommem[4598] <= 16'h0000;
rommem[4599] <= 16'h0000;
rommem[4600] <= 16'h0000;
rommem[4601] <= 16'h0000;
rommem[4602] <= 16'h0000;
rommem[4603] <= 16'h0000;
rommem[4604] <= 16'h0000;
rommem[4605] <= 16'h0000;
rommem[4606] <= 16'h0000;
rommem[4607] <= 16'h0000;
rommem[4608] <= 16'h0000;
rommem[4609] <= 16'h0000;
rommem[4610] <= 16'h0000;
rommem[4611] <= 16'h0000;
rommem[4612] <= 16'h0000;
rommem[4613] <= 16'h0000;
rommem[4614] <= 16'h0000;
rommem[4615] <= 16'h0000;
rommem[4616] <= 16'h0000;
rommem[4617] <= 16'h0000;
rommem[4618] <= 16'hFFFF;
rommem[4619] <= 16'hFFFF;
rommem[4620] <= 16'hFFFF;
rommem[4621] <= 16'hFFFF;
rommem[4622] <= 16'hFFFF;
rommem[4623] <= 16'hFFFF;
rommem[4624] <= 16'hFFFF;
rommem[4625] <= 16'hFFFF;
rommem[4626] <= 16'hFFFF;
rommem[4627] <= 16'hFFFF;
rommem[4628] <= 16'hFFFF;
rommem[4629] <= 16'hFFFF;
rommem[4630] <= 16'hFFFF;
rommem[4631] <= 16'hFFFF;
rommem[4632] <= 16'hFFFF;
rommem[4633] <= 16'hFFFF;
rommem[4634] <= 16'hFFFF;
rommem[4635] <= 16'hFFFF;
rommem[4636] <= 16'hFFFF;
rommem[4637] <= 16'hFFFF;
rommem[4638] <= 16'hFFFF;
rommem[4639] <= 16'hFFFF;
rommem[4640] <= 16'hFFFF;
rommem[4641] <= 16'hFFFF;
rommem[4642] <= 16'hFFFF;
rommem[4643] <= 16'hFFFF;
rommem[4644] <= 16'hFFFF;
rommem[4645] <= 16'hFFFF;
rommem[4646] <= 16'hFFFF;
rommem[4647] <= 16'hFFFF;
rommem[4648] <= 16'hFFFF;
rommem[4649] <= 16'hFFFF;
rommem[4650] <= 16'hFFFF;
rommem[4651] <= 16'hFFFF;
rommem[4652] <= 16'hFFFF;
rommem[4653] <= 16'hFFFF;
rommem[4654] <= 16'hFFFF;
rommem[4655] <= 16'hFFFF;
rommem[4656] <= 16'hFFFF;
rommem[4657] <= 16'hFFFF;
rommem[4658] <= 16'hFFFF;
rommem[4659] <= 16'hFFFF;
rommem[4660] <= 16'hFFFF;
rommem[4661] <= 16'hFFFF;
rommem[4662] <= 16'hFFFF;
rommem[4663] <= 16'hFFFF;
rommem[4664] <= 16'hFFFF;
rommem[4665] <= 16'hFFFF;
rommem[4666] <= 16'hFFFF;
rommem[4667] <= 16'hFFFF;
rommem[4668] <= 16'hFFFF;
rommem[4669] <= 16'hFFFF;
rommem[4670] <= 16'hFFFF;
rommem[4671] <= 16'hFFFF;
rommem[4672] <= 16'hFFFF;
rommem[4673] <= 16'hFFFF;
rommem[4674] <= 16'hFFFF;
rommem[4675] <= 16'hFFFF;
rommem[4676] <= 16'hFFFF;
rommem[4677] <= 16'hFFFF;
rommem[4678] <= 16'hFFFF;
rommem[4679] <= 16'hFFFF;
rommem[4680] <= 16'hFFFF;
rommem[4681] <= 16'hFFFF;
rommem[4682] <= 16'hFFFF;
rommem[4683] <= 16'hFFFF;
rommem[4684] <= 16'hFFFF;
rommem[4685] <= 16'hFFFF;
rommem[4686] <= 16'hFFFF;
rommem[4687] <= 16'hFFFF;
rommem[4688] <= 16'hFFFF;
rommem[4689] <= 16'hFFFF;
rommem[4690] <= 16'hFFFF;
rommem[4691] <= 16'hFFFF;
rommem[4692] <= 16'hFFFF;
rommem[4693] <= 16'hFFFF;
rommem[4694] <= 16'hFFFF;
rommem[4695] <= 16'hFFFF;
rommem[4696] <= 16'hFFFF;
rommem[4697] <= 16'hFFFF;
rommem[4698] <= 16'hFFFF;
rommem[4699] <= 16'hFFFF;
rommem[4700] <= 16'hFFFF;
rommem[4701] <= 16'hFFFF;
rommem[4702] <= 16'hFFFF;
rommem[4703] <= 16'hFFFF;
rommem[4704] <= 16'hFFFF;
rommem[4705] <= 16'hFFFF;
rommem[4706] <= 16'hFFFF;
rommem[4707] <= 16'hFFFF;
rommem[4708] <= 16'hFFFF;
rommem[4709] <= 16'hFFFF;
rommem[4710] <= 16'hFFFF;
rommem[4711] <= 16'hFFFF;
rommem[4712] <= 16'hFFFF;
rommem[4713] <= 16'hFFFF;
rommem[4714] <= 16'hFFFF;
rommem[4715] <= 16'hFFFF;
rommem[4716] <= 16'hFFFF;
rommem[4717] <= 16'hFFFF;
rommem[4718] <= 16'hFFFF;
rommem[4719] <= 16'hFFFF;
rommem[4720] <= 16'hFFFF;
rommem[4721] <= 16'hFFFF;
rommem[4722] <= 16'hFFFF;
rommem[4723] <= 16'hFFFF;
rommem[4724] <= 16'hFFFF;
rommem[4725] <= 16'hFFFF;
rommem[4726] <= 16'hFFFF;
rommem[4727] <= 16'hFFFF;
rommem[4728] <= 16'hFFFF;
rommem[4729] <= 16'hFFFF;
rommem[4730] <= 16'hFFFF;
rommem[4731] <= 16'hFFFF;
rommem[4732] <= 16'hFFFF;
rommem[4733] <= 16'hFFFF;
rommem[4734] <= 16'hFFFF;
rommem[4735] <= 16'hFFFF;
rommem[4736] <= 16'hFFFF;
rommem[4737] <= 16'hFFFF;
rommem[4738] <= 16'hFFFF;
rommem[4739] <= 16'hFFFF;
rommem[4740] <= 16'hFFFF;
rommem[4741] <= 16'hFFFF;
rommem[4742] <= 16'hFFFF;
rommem[4743] <= 16'hFFFF;
rommem[4744] <= 16'hFFFF;
rommem[4745] <= 16'hFFFF;
rommem[4746] <= 16'hFFFF;
rommem[4747] <= 16'hFFFF;
rommem[4748] <= 16'hFFFF;
rommem[4749] <= 16'hFFFF;
rommem[4750] <= 16'hFFFF;
rommem[4751] <= 16'hFFFF;
rommem[4752] <= 16'hFFFF;
rommem[4753] <= 16'hFFFF;
rommem[4754] <= 16'hFFFF;
rommem[4755] <= 16'hFFFF;
rommem[4756] <= 16'hFFFF;
rommem[4757] <= 16'hFFFF;
rommem[4758] <= 16'hFFFF;
rommem[4759] <= 16'hFFFF;
rommem[4760] <= 16'hFFFF;
rommem[4761] <= 16'hFFFF;
rommem[4762] <= 16'hFFFF;
rommem[4763] <= 16'hFFFF;
rommem[4764] <= 16'hFFFF;
rommem[4765] <= 16'hFFFF;
rommem[4766] <= 16'hFFFF;
rommem[4767] <= 16'hFFFF;
rommem[4768] <= 16'hFFFF;
rommem[4769] <= 16'hFFFF;
rommem[4770] <= 16'hFFFF;
rommem[4771] <= 16'hFFFF;
rommem[4772] <= 16'hFFFF;
rommem[4773] <= 16'hFFFF;
rommem[4774] <= 16'hFFFF;
rommem[4775] <= 16'hFFFF;
rommem[4776] <= 16'hFFFF;
rommem[4777] <= 16'hFFFF;
rommem[4778] <= 16'hFFFF;
rommem[4779] <= 16'hFFFF;
rommem[4780] <= 16'hFFFF;
rommem[4781] <= 16'hFFFF;
rommem[4782] <= 16'hFFFF;
rommem[4783] <= 16'hFFFF;
rommem[4784] <= 16'hFFFF;
rommem[4785] <= 16'hFFFF;
rommem[4786] <= 16'hFFFF;
rommem[4787] <= 16'hFFFF;
rommem[4788] <= 16'hFFFF;
rommem[4789] <= 16'hFFFF;
rommem[4790] <= 16'hFFFF;
rommem[4791] <= 16'hFFFF;
rommem[4792] <= 16'hFFFF;
rommem[4793] <= 16'hFFFF;
rommem[4794] <= 16'hFFFF;
rommem[4795] <= 16'hFFFF;
rommem[4796] <= 16'hFFFF;
rommem[4797] <= 16'hFFFF;
rommem[4798] <= 16'hFFFF;
rommem[4799] <= 16'hFFFF;
rommem[4800] <= 16'hFFFF;
rommem[4801] <= 16'hFFFF;
rommem[4802] <= 16'hFFFF;
rommem[4803] <= 16'hFFFF;
rommem[4804] <= 16'hFFFF;
rommem[4805] <= 16'hFFFF;
rommem[4806] <= 16'hFFFF;
rommem[4807] <= 16'hFFFF;
rommem[4808] <= 16'hFFFF;
rommem[4809] <= 16'hFFFF;
rommem[4810] <= 16'hFFFF;
rommem[4811] <= 16'hFFFF;
rommem[4812] <= 16'hFFFF;
rommem[4813] <= 16'hFFFF;
rommem[4814] <= 16'hFFFF;
rommem[4815] <= 16'hFFFF;
rommem[4816] <= 16'hFFFF;
rommem[4817] <= 16'hFFFF;
rommem[4818] <= 16'hFFFF;
rommem[4819] <= 16'hFFFF;
rommem[4820] <= 16'hFFFF;
rommem[4821] <= 16'hFFFF;
rommem[4822] <= 16'hFFFF;
rommem[4823] <= 16'hFFFF;
rommem[4824] <= 16'hFFFF;
rommem[4825] <= 16'hFFFF;
rommem[4826] <= 16'hFFFF;
rommem[4827] <= 16'hFFFF;
rommem[4828] <= 16'hFFFF;
rommem[4829] <= 16'hFFFF;
rommem[4830] <= 16'hFFFF;
rommem[4831] <= 16'hFFFF;
rommem[4832] <= 16'hFFFF;
rommem[4833] <= 16'hFFFF;
rommem[4834] <= 16'hFFFF;
rommem[4835] <= 16'hFFFF;
rommem[4836] <= 16'hFFFF;
rommem[4837] <= 16'hFFFF;
rommem[4838] <= 16'hFFFF;
rommem[4839] <= 16'hFFFF;
rommem[4840] <= 16'hFFFF;
rommem[4841] <= 16'hFFFF;
rommem[4842] <= 16'hFFFF;
rommem[4843] <= 16'hFFFF;
rommem[4844] <= 16'hFFFF;
rommem[4845] <= 16'hFFFF;
rommem[4846] <= 16'hFFFF;
rommem[4847] <= 16'hFFFF;
rommem[4848] <= 16'hFFFF;
rommem[4849] <= 16'hFFFF;
rommem[4850] <= 16'hFFFF;
rommem[4851] <= 16'hFFFF;
rommem[4852] <= 16'hFFFF;
rommem[4853] <= 16'hFFFF;
rommem[4854] <= 16'hFFFF;
rommem[4855] <= 16'hFFFF;
rommem[4856] <= 16'hFFFF;
rommem[4857] <= 16'hFFFF;
rommem[4858] <= 16'hFFFF;
rommem[4859] <= 16'hFFFF;
rommem[4860] <= 16'hFFFF;
rommem[4861] <= 16'hFFFF;
rommem[4862] <= 16'hFFFF;
rommem[4863] <= 16'hFFFF;
rommem[4864] <= 16'hFFFF;
rommem[4865] <= 16'hFFFF;
rommem[4866] <= 16'hFFFF;
rommem[4867] <= 16'hFFFF;
rommem[4868] <= 16'hFFFF;
rommem[4869] <= 16'hFFFF;
rommem[4870] <= 16'hFFFF;
rommem[4871] <= 16'hFFFF;
rommem[4872] <= 16'hFFFF;
rommem[4873] <= 16'hFFFF;
rommem[4874] <= 16'hFFFF;
rommem[4875] <= 16'hFFFF;
rommem[4876] <= 16'hFFFF;
rommem[4877] <= 16'hFFFF;
rommem[4878] <= 16'hFFFF;
rommem[4879] <= 16'hFFFF;
rommem[4880] <= 16'hFFFF;
rommem[4881] <= 16'hFFFF;
rommem[4882] <= 16'hFFFF;
rommem[4883] <= 16'hFFFF;
rommem[4884] <= 16'hFFFF;
rommem[4885] <= 16'hFFFF;
rommem[4886] <= 16'hFFFF;
rommem[4887] <= 16'hFFFF;
rommem[4888] <= 16'hFFFF;
rommem[4889] <= 16'hFFFF;
rommem[4890] <= 16'hFFFF;
rommem[4891] <= 16'hFFFF;
rommem[4892] <= 16'hFFFF;
rommem[4893] <= 16'hFFFF;
rommem[4894] <= 16'hFFFF;
rommem[4895] <= 16'hFFFF;
rommem[4896] <= 16'hFFFF;
rommem[4897] <= 16'hFFFF;
rommem[4898] <= 16'hFFFF;
rommem[4899] <= 16'hFFFF;
rommem[4900] <= 16'hFFFF;
rommem[4901] <= 16'hFFFF;
rommem[4902] <= 16'hFFFF;
rommem[4903] <= 16'hFFFF;
rommem[4904] <= 16'hFFFF;
rommem[4905] <= 16'hFFFF;
rommem[4906] <= 16'hFFFF;
rommem[4907] <= 16'hFFFF;
rommem[4908] <= 16'hFFFF;
rommem[4909] <= 16'hFFFF;
rommem[4910] <= 16'hFFFF;
rommem[4911] <= 16'hFFFF;
rommem[4912] <= 16'hFFFF;
rommem[4913] <= 16'hFFFF;
rommem[4914] <= 16'hFFFF;
rommem[4915] <= 16'hFFFF;
rommem[4916] <= 16'hFFFF;
rommem[4917] <= 16'hFFFF;
rommem[4918] <= 16'hFFFF;
rommem[4919] <= 16'hFFFF;
rommem[4920] <= 16'hFFFF;
rommem[4921] <= 16'hFFFF;
rommem[4922] <= 16'hFFFF;
rommem[4923] <= 16'hFFFF;
rommem[4924] <= 16'hFFFF;
rommem[4925] <= 16'hFFFF;
rommem[4926] <= 16'hFFFF;
rommem[4927] <= 16'hFFFF;
rommem[4928] <= 16'hFFFF;
rommem[4929] <= 16'hFFFF;
rommem[4930] <= 16'hFFFF;
rommem[4931] <= 16'hFFFF;
rommem[4932] <= 16'hFFFF;
rommem[4933] <= 16'hFFFF;
rommem[4934] <= 16'hFFFF;
rommem[4935] <= 16'hFFFF;
rommem[4936] <= 16'hFFFF;
rommem[4937] <= 16'hFFFF;
rommem[4938] <= 16'hFFFF;
rommem[4939] <= 16'hFFFF;
rommem[4940] <= 16'hFFFF;
rommem[4941] <= 16'hFFFF;
rommem[4942] <= 16'hFFFF;
rommem[4943] <= 16'hFFFF;
rommem[4944] <= 16'hFFFF;
rommem[4945] <= 16'hFFFF;
rommem[4946] <= 16'hFFFF;
rommem[4947] <= 16'hFFFF;
rommem[4948] <= 16'hFFFF;
rommem[4949] <= 16'hFFFF;
rommem[4950] <= 16'hFFFF;
rommem[4951] <= 16'hFFFF;
rommem[4952] <= 16'hFFFF;
rommem[4953] <= 16'hFFFF;
rommem[4954] <= 16'hFFFF;
rommem[4955] <= 16'hFFFF;
rommem[4956] <= 16'hFFFF;
rommem[4957] <= 16'hFFFF;
rommem[4958] <= 16'hFFFF;
rommem[4959] <= 16'hFFFF;
rommem[4960] <= 16'hFFFF;
rommem[4961] <= 16'hFFFF;
rommem[4962] <= 16'hFFFF;
rommem[4963] <= 16'hFFFF;
rommem[4964] <= 16'hFFFF;
rommem[4965] <= 16'hFFFF;
rommem[4966] <= 16'hFFFF;
rommem[4967] <= 16'hFFFF;
rommem[4968] <= 16'hFFFF;
rommem[4969] <= 16'hFFFF;
rommem[4970] <= 16'hFFFF;
rommem[4971] <= 16'hFFFF;
rommem[4972] <= 16'hFFFF;
rommem[4973] <= 16'hFFFF;
rommem[4974] <= 16'hFFFF;
rommem[4975] <= 16'hFFFF;
rommem[4976] <= 16'hFFFF;
rommem[4977] <= 16'hFFFF;
rommem[4978] <= 16'hFFFF;
rommem[4979] <= 16'hFFFF;
rommem[4980] <= 16'hFFFF;
rommem[4981] <= 16'hFFFF;
rommem[4982] <= 16'hFFFF;
rommem[4983] <= 16'hFFFF;
rommem[4984] <= 16'hFFFF;
rommem[4985] <= 16'hFFFF;
rommem[4986] <= 16'hFFFF;
rommem[4987] <= 16'hFFFF;
rommem[4988] <= 16'hFFFF;
rommem[4989] <= 16'hFFFF;
rommem[4990] <= 16'hFFFF;
rommem[4991] <= 16'hFFFF;
rommem[4992] <= 16'hFFFF;
rommem[4993] <= 16'hFFFF;
rommem[4994] <= 16'hFFFF;
rommem[4995] <= 16'hFFFF;
rommem[4996] <= 16'hFFFF;
rommem[4997] <= 16'hFFFF;
rommem[4998] <= 16'hFFFF;
rommem[4999] <= 16'hFFFF;
rommem[5000] <= 16'hFFFF;
rommem[5001] <= 16'hFFFF;
rommem[5002] <= 16'hFFFF;
rommem[5003] <= 16'hFFFF;
rommem[5004] <= 16'hFFFF;
rommem[5005] <= 16'hFFFF;
rommem[5006] <= 16'hFFFF;
rommem[5007] <= 16'hFFFF;
rommem[5008] <= 16'hFFFF;
rommem[5009] <= 16'hFFFF;
rommem[5010] <= 16'hFFFF;
rommem[5011] <= 16'hFFFF;
rommem[5012] <= 16'hFFFF;
rommem[5013] <= 16'hFFFF;
rommem[5014] <= 16'hFFFF;
rommem[5015] <= 16'hFFFF;
rommem[5016] <= 16'hFFFF;
rommem[5017] <= 16'hFFFF;
rommem[5018] <= 16'hFFFF;
rommem[5019] <= 16'hFFFF;
rommem[5020] <= 16'hFFFF;
rommem[5021] <= 16'hFFFF;
rommem[5022] <= 16'hFFFF;
rommem[5023] <= 16'hFFFF;
rommem[5024] <= 16'hFFFF;
rommem[5025] <= 16'hFFFF;
rommem[5026] <= 16'hFFFF;
rommem[5027] <= 16'hFFFF;
rommem[5028] <= 16'hFFFF;
rommem[5029] <= 16'hFFFF;
rommem[5030] <= 16'hFFFF;
rommem[5031] <= 16'hFFFF;
rommem[5032] <= 16'hFFFF;
rommem[5033] <= 16'hFFFF;
rommem[5034] <= 16'hFFFF;
rommem[5035] <= 16'hFFFF;
rommem[5036] <= 16'hFFFF;
rommem[5037] <= 16'hFFFF;
rommem[5038] <= 16'hFFFF;
rommem[5039] <= 16'hFFFF;
rommem[5040] <= 16'hFFFF;
rommem[5041] <= 16'hFFFF;
rommem[5042] <= 16'hFFFF;
rommem[5043] <= 16'hFFFF;
rommem[5044] <= 16'hFFFF;
rommem[5045] <= 16'hFFFF;
rommem[5046] <= 16'hFFFF;
rommem[5047] <= 16'hFFFF;
rommem[5048] <= 16'hFFFF;
rommem[5049] <= 16'hFFFF;
rommem[5050] <= 16'hFFFF;
rommem[5051] <= 16'hFFFF;
rommem[5052] <= 16'hFFFF;
rommem[5053] <= 16'hFFFF;
rommem[5054] <= 16'hFFFF;
rommem[5055] <= 16'hFFFF;
rommem[5056] <= 16'hFFFF;
rommem[5057] <= 16'hFFFF;
rommem[5058] <= 16'hFFFF;
rommem[5059] <= 16'hFFFF;
rommem[5060] <= 16'hFFFF;
rommem[5061] <= 16'hFFFF;
rommem[5062] <= 16'hFFFF;
rommem[5063] <= 16'hFFFF;
rommem[5064] <= 16'hFFFF;
rommem[5065] <= 16'hFFFF;
rommem[5066] <= 16'hFFFF;
rommem[5067] <= 16'hFFFF;
rommem[5068] <= 16'hFFFF;
rommem[5069] <= 16'hFFFF;
rommem[5070] <= 16'hFFFF;
rommem[5071] <= 16'hFFFF;
rommem[5072] <= 16'hFFFF;
rommem[5073] <= 16'hFFFF;
rommem[5074] <= 16'hFFFF;
rommem[5075] <= 16'hFFFF;
rommem[5076] <= 16'hFFFF;
rommem[5077] <= 16'hFFFF;
rommem[5078] <= 16'hFFFF;
rommem[5079] <= 16'hFFFF;
rommem[5080] <= 16'hFFFF;
rommem[5081] <= 16'hFFFF;
rommem[5082] <= 16'hFFFF;
rommem[5083] <= 16'hFFFF;
rommem[5084] <= 16'hFFFF;
rommem[5085] <= 16'hFFFF;
rommem[5086] <= 16'hFFFF;
rommem[5087] <= 16'hFFFF;
rommem[5088] <= 16'hFFFF;
rommem[5089] <= 16'hFFFF;
rommem[5090] <= 16'hFFFF;
rommem[5091] <= 16'hFFFF;
rommem[5092] <= 16'hFFFF;
rommem[5093] <= 16'hFFFF;
rommem[5094] <= 16'hFFFF;
rommem[5095] <= 16'hFFFF;
rommem[5096] <= 16'hFFFF;
rommem[5097] <= 16'hFFFF;
rommem[5098] <= 16'hFFFF;
rommem[5099] <= 16'hFFFF;
rommem[5100] <= 16'hFFFF;
rommem[5101] <= 16'hFFFF;
rommem[5102] <= 16'hFFFF;
rommem[5103] <= 16'hFFFF;
rommem[5104] <= 16'hFFFF;
rommem[5105] <= 16'hFFFF;
rommem[5106] <= 16'hFFFF;
rommem[5107] <= 16'hFFFF;
rommem[5108] <= 16'hFFFF;
rommem[5109] <= 16'hFFFF;
rommem[5110] <= 16'hFFFF;
rommem[5111] <= 16'hFFFF;
rommem[5112] <= 16'hFFFF;
rommem[5113] <= 16'hFFFF;
rommem[5114] <= 16'hFFFF;
rommem[5115] <= 16'hFFFF;
rommem[5116] <= 16'hFFFF;
rommem[5117] <= 16'hFFFF;
rommem[5118] <= 16'hFFFF;
rommem[5119] <= 16'hFFFF;
rommem[5120] <= 16'hFFFF;
rommem[5121] <= 16'hFFFF;
rommem[5122] <= 16'hFFFF;
rommem[5123] <= 16'hFFFF;
rommem[5124] <= 16'hFFFF;
rommem[5125] <= 16'hFFFF;
rommem[5126] <= 16'hFFFF;
rommem[5127] <= 16'hFFFF;
rommem[5128] <= 16'hFFFF;
rommem[5129] <= 16'hFFFF;
rommem[5130] <= 16'hFFFF;
rommem[5131] <= 16'hFFFF;
rommem[5132] <= 16'hFFFF;
rommem[5133] <= 16'hFFFF;
rommem[5134] <= 16'hFFFF;
rommem[5135] <= 16'hFFFF;
rommem[5136] <= 16'hFFFF;
rommem[5137] <= 16'hFFFF;
rommem[5138] <= 16'hFFFF;
rommem[5139] <= 16'hFFFF;
rommem[5140] <= 16'hFFFF;
rommem[5141] <= 16'hFFFF;
rommem[5142] <= 16'hFFFF;
rommem[5143] <= 16'hFFFF;
rommem[5144] <= 16'hFFFF;
rommem[5145] <= 16'hFFFF;
rommem[5146] <= 16'hFFFF;
rommem[5147] <= 16'hFFFF;
rommem[5148] <= 16'hFFFF;
rommem[5149] <= 16'hFFFF;
rommem[5150] <= 16'hFFFF;
rommem[5151] <= 16'hFFFF;
rommem[5152] <= 16'hFFFF;
rommem[5153] <= 16'hFFFF;
rommem[5154] <= 16'hFFFF;
rommem[5155] <= 16'hFFFF;
rommem[5156] <= 16'hFFFF;
rommem[5157] <= 16'hFFFF;
rommem[5158] <= 16'hFFFF;
rommem[5159] <= 16'hFFFF;
rommem[5160] <= 16'hFFFF;
rommem[5161] <= 16'hFFFF;
rommem[5162] <= 16'hFFFF;
rommem[5163] <= 16'hFFFF;
rommem[5164] <= 16'hFFFF;
rommem[5165] <= 16'hFFFF;
rommem[5166] <= 16'hFFFF;
rommem[5167] <= 16'hFFFF;
rommem[5168] <= 16'hFFFF;
rommem[5169] <= 16'hFFFF;
rommem[5170] <= 16'hFFFF;
rommem[5171] <= 16'hFFFF;
rommem[5172] <= 16'hFFFF;
rommem[5173] <= 16'hFFFF;
rommem[5174] <= 16'hFFFF;
rommem[5175] <= 16'hFFFF;
rommem[5176] <= 16'hFFFF;
rommem[5177] <= 16'hFFFF;
rommem[5178] <= 16'hFFFF;
rommem[5179] <= 16'hFFFF;
rommem[5180] <= 16'hFFFF;
rommem[5181] <= 16'hFFFF;
rommem[5182] <= 16'hFFFF;
rommem[5183] <= 16'hFFFF;
rommem[5184] <= 16'hFFFF;
rommem[5185] <= 16'hFFFF;
rommem[5186] <= 16'hFFFF;
rommem[5187] <= 16'hFFFF;
rommem[5188] <= 16'hFFFF;
rommem[5189] <= 16'hFFFF;
rommem[5190] <= 16'hFFFF;
rommem[5191] <= 16'hFFFF;
rommem[5192] <= 16'hFFFF;
rommem[5193] <= 16'hFFFF;
rommem[5194] <= 16'hFFFF;
rommem[5195] <= 16'hFFFF;
rommem[5196] <= 16'hFFFF;
rommem[5197] <= 16'hFFFF;
rommem[5198] <= 16'hFFFF;
rommem[5199] <= 16'hFFFF;
rommem[5200] <= 16'hFFFF;
rommem[5201] <= 16'hFFFF;
rommem[5202] <= 16'hFFFF;
rommem[5203] <= 16'hFFFF;
rommem[5204] <= 16'hFFFF;
rommem[5205] <= 16'hFFFF;
rommem[5206] <= 16'hFFFF;
rommem[5207] <= 16'hFFFF;
rommem[5208] <= 16'hFFFF;
rommem[5209] <= 16'hFFFF;
rommem[5210] <= 16'hFFFF;
rommem[5211] <= 16'hFFFF;
rommem[5212] <= 16'hFFFF;
rommem[5213] <= 16'hFFFF;
rommem[5214] <= 16'hFFFF;
rommem[5215] <= 16'hFFFF;
rommem[5216] <= 16'hFFFF;
rommem[5217] <= 16'hFFFF;
rommem[5218] <= 16'hFFFF;
rommem[5219] <= 16'hFFFF;
rommem[5220] <= 16'hFFFF;
rommem[5221] <= 16'hFFFF;
rommem[5222] <= 16'hFFFF;
rommem[5223] <= 16'hFFFF;
rommem[5224] <= 16'hFFFF;
rommem[5225] <= 16'hFFFF;
rommem[5226] <= 16'hFFFF;
rommem[5227] <= 16'hFFFF;
rommem[5228] <= 16'hFFFF;
rommem[5229] <= 16'hFFFF;
rommem[5230] <= 16'hFFFF;
rommem[5231] <= 16'hFFFF;
rommem[5232] <= 16'hFFFF;
rommem[5233] <= 16'hFFFF;
rommem[5234] <= 16'hFFFF;
rommem[5235] <= 16'hFFFF;
rommem[5236] <= 16'hFFFF;
rommem[5237] <= 16'hFFFF;
rommem[5238] <= 16'hFFFF;
rommem[5239] <= 16'hFFFF;
rommem[5240] <= 16'hFFFF;
rommem[5241] <= 16'hFFFF;
rommem[5242] <= 16'hFFFF;
rommem[5243] <= 16'hFFFF;
rommem[5244] <= 16'hFFFF;
rommem[5245] <= 16'hFFFF;
rommem[5246] <= 16'hFFFF;
rommem[5247] <= 16'hFFFF;
rommem[5248] <= 16'hFFFF;
rommem[5249] <= 16'hFFFF;
rommem[5250] <= 16'hFFFF;
rommem[5251] <= 16'hFFFF;
rommem[5252] <= 16'hFFFF;
rommem[5253] <= 16'hFFFF;
rommem[5254] <= 16'hFFFF;
rommem[5255] <= 16'hFFFF;
rommem[5256] <= 16'hFFFF;
rommem[5257] <= 16'hFFFF;
rommem[5258] <= 16'hFFFF;
rommem[5259] <= 16'hFFFF;
rommem[5260] <= 16'hFFFF;
rommem[5261] <= 16'hFFFF;
rommem[5262] <= 16'hFFFF;
rommem[5263] <= 16'hFFFF;
rommem[5264] <= 16'hFFFF;
rommem[5265] <= 16'hFFFF;
rommem[5266] <= 16'hFFFF;
rommem[5267] <= 16'hFFFF;
rommem[5268] <= 16'hFFFF;
rommem[5269] <= 16'hFFFF;
rommem[5270] <= 16'hFFFF;
rommem[5271] <= 16'hFFFF;
rommem[5272] <= 16'hFFFF;
rommem[5273] <= 16'hFFFF;
rommem[5274] <= 16'hFFFF;
rommem[5275] <= 16'hFFFF;
rommem[5276] <= 16'hFFFF;
rommem[5277] <= 16'hFFFF;
rommem[5278] <= 16'hFFFF;
rommem[5279] <= 16'hFFFF;
rommem[5280] <= 16'hFFFF;
rommem[5281] <= 16'hFFFF;
rommem[5282] <= 16'hFFFF;
rommem[5283] <= 16'hFFFF;
rommem[5284] <= 16'hFFFF;
rommem[5285] <= 16'hFFFF;
rommem[5286] <= 16'hFFFF;
rommem[5287] <= 16'hFFFF;
rommem[5288] <= 16'hFFFF;
rommem[5289] <= 16'hFFFF;
rommem[5290] <= 16'hFFFF;
rommem[5291] <= 16'hFFFF;
rommem[5292] <= 16'hFFFF;
rommem[5293] <= 16'hFFFF;
rommem[5294] <= 16'hFFFF;
rommem[5295] <= 16'hFFFF;
rommem[5296] <= 16'hFFFF;
rommem[5297] <= 16'hFFFF;
rommem[5298] <= 16'hFFFF;
rommem[5299] <= 16'hFFFF;
rommem[5300] <= 16'hFFFF;
rommem[5301] <= 16'hFFFF;
rommem[5302] <= 16'hFFFF;
rommem[5303] <= 16'hFFFF;
rommem[5304] <= 16'hFFFF;
rommem[5305] <= 16'hFFFF;
rommem[5306] <= 16'hFFFF;
rommem[5307] <= 16'hFFFF;
rommem[5308] <= 16'hFFFF;
rommem[5309] <= 16'hFFFF;
rommem[5310] <= 16'hFFFF;
rommem[5311] <= 16'hFFFF;
rommem[5312] <= 16'hFFFF;
rommem[5313] <= 16'hFFFF;
rommem[5314] <= 16'hFFFF;
rommem[5315] <= 16'hFFFF;
rommem[5316] <= 16'hFFFF;
rommem[5317] <= 16'hFFFF;
rommem[5318] <= 16'hFFFF;
rommem[5319] <= 16'hFFFF;
rommem[5320] <= 16'hFFFF;
rommem[5321] <= 16'hFFFF;
rommem[5322] <= 16'hFFFF;
rommem[5323] <= 16'hFFFF;
rommem[5324] <= 16'hFFFF;
rommem[5325] <= 16'hFFFF;
rommem[5326] <= 16'hFFFF;
rommem[5327] <= 16'hFFFF;
rommem[5328] <= 16'hFFFF;
rommem[5329] <= 16'hFFFF;
rommem[5330] <= 16'hFFFF;
rommem[5331] <= 16'hFFFF;
rommem[5332] <= 16'hFFFF;
rommem[5333] <= 16'hFFFF;
rommem[5334] <= 16'hFFFF;
rommem[5335] <= 16'hFFFF;
rommem[5336] <= 16'hFFFF;
rommem[5337] <= 16'hFFFF;
rommem[5338] <= 16'hFFFF;
rommem[5339] <= 16'hFFFF;
rommem[5340] <= 16'hFFFF;
rommem[5341] <= 16'hFFFF;
rommem[5342] <= 16'hFFFF;
rommem[5343] <= 16'hFFFF;
rommem[5344] <= 16'hFFFF;
rommem[5345] <= 16'hFFFF;
rommem[5346] <= 16'hFFFF;
rommem[5347] <= 16'hFFFF;
rommem[5348] <= 16'hFFFF;
rommem[5349] <= 16'hFFFF;
rommem[5350] <= 16'hFFFF;
rommem[5351] <= 16'hFFFF;
rommem[5352] <= 16'hFFFF;
rommem[5353] <= 16'hFFFF;
rommem[5354] <= 16'hFFFF;
rommem[5355] <= 16'hFFFF;
rommem[5356] <= 16'hFFFF;
rommem[5357] <= 16'hFFFF;
rommem[5358] <= 16'hFFFF;
rommem[5359] <= 16'hFFFF;
rommem[5360] <= 16'hFFFF;
rommem[5361] <= 16'hFFFF;
rommem[5362] <= 16'hFFFF;
rommem[5363] <= 16'hFFFF;
rommem[5364] <= 16'hFFFF;
rommem[5365] <= 16'hFFFF;
rommem[5366] <= 16'hFFFF;
rommem[5367] <= 16'hFFFF;
rommem[5368] <= 16'hFFFF;
rommem[5369] <= 16'hFFFF;
rommem[5370] <= 16'hFFFF;
rommem[5371] <= 16'hFFFF;
rommem[5372] <= 16'hFFFF;
rommem[5373] <= 16'hFFFF;
rommem[5374] <= 16'hFFFF;
rommem[5375] <= 16'hFFFF;
rommem[5376] <= 16'hFFFF;
rommem[5377] <= 16'hFFFF;
rommem[5378] <= 16'hFFFF;
rommem[5379] <= 16'hFFFF;
rommem[5380] <= 16'hFFFF;
rommem[5381] <= 16'hFFFF;
rommem[5382] <= 16'hFFFF;
rommem[5383] <= 16'hFFFF;
rommem[5384] <= 16'hFFFF;
rommem[5385] <= 16'hFFFF;
rommem[5386] <= 16'hFFFF;
rommem[5387] <= 16'hFFFF;
rommem[5388] <= 16'hFFFF;
rommem[5389] <= 16'hFFFF;
rommem[5390] <= 16'hFFFF;
rommem[5391] <= 16'hFFFF;
rommem[5392] <= 16'hFFFF;
rommem[5393] <= 16'hFFFF;
rommem[5394] <= 16'hFFFF;
rommem[5395] <= 16'hFFFF;
rommem[5396] <= 16'hFFFF;
rommem[5397] <= 16'hFFFF;
rommem[5398] <= 16'hFFFF;
rommem[5399] <= 16'hFFFF;
rommem[5400] <= 16'hFFFF;
rommem[5401] <= 16'hFFFF;
rommem[5402] <= 16'hFFFF;
rommem[5403] <= 16'hFFFF;
rommem[5404] <= 16'hFFFF;
rommem[5405] <= 16'hFFFF;
rommem[5406] <= 16'hFFFF;
rommem[5407] <= 16'hFFFF;
rommem[5408] <= 16'hFFFF;
rommem[5409] <= 16'hFFFF;
rommem[5410] <= 16'hFFFF;
rommem[5411] <= 16'hFFFF;
rommem[5412] <= 16'hFFFF;
rommem[5413] <= 16'hFFFF;
rommem[5414] <= 16'hFFFF;
rommem[5415] <= 16'hFFFF;
rommem[5416] <= 16'hFFFF;
rommem[5417] <= 16'hFFFF;
rommem[5418] <= 16'hFFFF;
rommem[5419] <= 16'hFFFF;
rommem[5420] <= 16'hFFFF;
rommem[5421] <= 16'hFFFF;
rommem[5422] <= 16'hFFFF;
rommem[5423] <= 16'hFFFF;
rommem[5424] <= 16'hFFFF;
rommem[5425] <= 16'hFFFF;
rommem[5426] <= 16'hFFFF;
rommem[5427] <= 16'hFFFF;
rommem[5428] <= 16'hFFFF;
rommem[5429] <= 16'hFFFF;
rommem[5430] <= 16'hFFFF;
rommem[5431] <= 16'hFFFF;
rommem[5432] <= 16'hFFFF;
rommem[5433] <= 16'hFFFF;
rommem[5434] <= 16'hFFFF;
rommem[5435] <= 16'hFFFF;
rommem[5436] <= 16'hFFFF;
rommem[5437] <= 16'hFFFF;
rommem[5438] <= 16'hFFFF;
rommem[5439] <= 16'hFFFF;
rommem[5440] <= 16'hFFFF;
rommem[5441] <= 16'hFFFF;
rommem[5442] <= 16'hFFFF;
rommem[5443] <= 16'hFFFF;
rommem[5444] <= 16'hFFFF;
rommem[5445] <= 16'hFFFF;
rommem[5446] <= 16'hFFFF;
rommem[5447] <= 16'hFFFF;
rommem[5448] <= 16'hFFFF;
rommem[5449] <= 16'hFFFF;
rommem[5450] <= 16'hFFFF;
rommem[5451] <= 16'hFFFF;
rommem[5452] <= 16'hFFFF;
rommem[5453] <= 16'hFFFF;
rommem[5454] <= 16'hFFFF;
rommem[5455] <= 16'hFFFF;
rommem[5456] <= 16'hFFFF;
rommem[5457] <= 16'hFFFF;
rommem[5458] <= 16'hFFFF;
rommem[5459] <= 16'hFFFF;
rommem[5460] <= 16'hFFFF;
rommem[5461] <= 16'hFFFF;
rommem[5462] <= 16'hFFFF;
rommem[5463] <= 16'hFFFF;
rommem[5464] <= 16'hFFFF;
rommem[5465] <= 16'hFFFF;
rommem[5466] <= 16'hFFFF;
rommem[5467] <= 16'hFFFF;
rommem[5468] <= 16'hFFFF;
rommem[5469] <= 16'hFFFF;
rommem[5470] <= 16'hFFFF;
rommem[5471] <= 16'hFFFF;
rommem[5472] <= 16'hFFFF;
rommem[5473] <= 16'hFFFF;
rommem[5474] <= 16'hFFFF;
rommem[5475] <= 16'hFFFF;
rommem[5476] <= 16'hFFFF;
rommem[5477] <= 16'hFFFF;
rommem[5478] <= 16'hFFFF;
rommem[5479] <= 16'hFFFF;
rommem[5480] <= 16'hFFFF;
rommem[5481] <= 16'hFFFF;
rommem[5482] <= 16'hFFFF;
rommem[5483] <= 16'hFFFF;
rommem[5484] <= 16'hFFFF;
rommem[5485] <= 16'hFFFF;
rommem[5486] <= 16'hFFFF;
rommem[5487] <= 16'hFFFF;
rommem[5488] <= 16'hFFFF;
rommem[5489] <= 16'hFFFF;
rommem[5490] <= 16'hFFFF;
rommem[5491] <= 16'hFFFF;
rommem[5492] <= 16'hFFFF;
rommem[5493] <= 16'hFFFF;
rommem[5494] <= 16'hFFFF;
rommem[5495] <= 16'hFFFF;
rommem[5496] <= 16'hFFFF;
rommem[5497] <= 16'hFFFF;
rommem[5498] <= 16'hFFFF;
rommem[5499] <= 16'hFFFF;
rommem[5500] <= 16'hFFFF;
rommem[5501] <= 16'hFFFF;
rommem[5502] <= 16'hFFFF;
rommem[5503] <= 16'hFFFF;
rommem[5504] <= 16'hFFFF;
rommem[5505] <= 16'hFFFF;
rommem[5506] <= 16'hFFFF;
rommem[5507] <= 16'hFFFF;
rommem[5508] <= 16'hFFFF;
rommem[5509] <= 16'hFFFF;
rommem[5510] <= 16'hFFFF;
rommem[5511] <= 16'hFFFF;
rommem[5512] <= 16'hFFFF;
rommem[5513] <= 16'hFFFF;
rommem[5514] <= 16'hFFFF;
rommem[5515] <= 16'hFFFF;
rommem[5516] <= 16'hFFFF;
rommem[5517] <= 16'hFFFF;
rommem[5518] <= 16'hFFFF;
rommem[5519] <= 16'hFFFF;
rommem[5520] <= 16'hFFFF;
rommem[5521] <= 16'hFFFF;
rommem[5522] <= 16'hFFFF;
rommem[5523] <= 16'hFFFF;
rommem[5524] <= 16'hFFFF;
rommem[5525] <= 16'hFFFF;
rommem[5526] <= 16'hFFFF;
rommem[5527] <= 16'hFFFF;
rommem[5528] <= 16'hFFFF;
rommem[5529] <= 16'hFFFF;
rommem[5530] <= 16'hFFFF;
rommem[5531] <= 16'hFFFF;
rommem[5532] <= 16'hFFFF;
rommem[5533] <= 16'hFFFF;
rommem[5534] <= 16'hFFFF;
rommem[5535] <= 16'hFFFF;
rommem[5536] <= 16'hFFFF;
rommem[5537] <= 16'hFFFF;
rommem[5538] <= 16'hFFFF;
rommem[5539] <= 16'hFFFF;
rommem[5540] <= 16'hFFFF;
rommem[5541] <= 16'hFFFF;
rommem[5542] <= 16'hFFFF;
rommem[5543] <= 16'hFFFF;
rommem[5544] <= 16'hFFFF;
rommem[5545] <= 16'hFFFF;
rommem[5546] <= 16'hFFFF;
rommem[5547] <= 16'hFFFF;
rommem[5548] <= 16'hFFFF;
rommem[5549] <= 16'hFFFF;
rommem[5550] <= 16'hFFFF;
rommem[5551] <= 16'hFFFF;
rommem[5552] <= 16'hFFFF;
rommem[5553] <= 16'hFFFF;
rommem[5554] <= 16'hFFFF;
rommem[5555] <= 16'hFFFF;
rommem[5556] <= 16'hFFFF;
rommem[5557] <= 16'hFFFF;
rommem[5558] <= 16'hFFFF;
rommem[5559] <= 16'hFFFF;
rommem[5560] <= 16'hFFFF;
rommem[5561] <= 16'hFFFF;
rommem[5562] <= 16'hFFFF;
rommem[5563] <= 16'hFFFF;
rommem[5564] <= 16'hFFFF;
rommem[5565] <= 16'hFFFF;
rommem[5566] <= 16'hFFFF;
rommem[5567] <= 16'hFFFF;
rommem[5568] <= 16'hFFFF;
rommem[5569] <= 16'hFFFF;
rommem[5570] <= 16'hFFFF;
rommem[5571] <= 16'hFFFF;
rommem[5572] <= 16'hFFFF;
rommem[5573] <= 16'hFFFF;
rommem[5574] <= 16'hFFFF;
rommem[5575] <= 16'hFFFF;
rommem[5576] <= 16'hFFFF;
rommem[5577] <= 16'hFFFF;
rommem[5578] <= 16'hFFFF;
rommem[5579] <= 16'hFFFF;
rommem[5580] <= 16'hFFFF;
rommem[5581] <= 16'hFFFF;
rommem[5582] <= 16'hFFFF;
rommem[5583] <= 16'hFFFF;
rommem[5584] <= 16'hFFFF;
rommem[5585] <= 16'hFFFF;
rommem[5586] <= 16'hFFFF;
rommem[5587] <= 16'hFFFF;
rommem[5588] <= 16'hFFFF;
rommem[5589] <= 16'hFFFF;
rommem[5590] <= 16'hFFFF;
rommem[5591] <= 16'hFFFF;
rommem[5592] <= 16'hFFFF;
rommem[5593] <= 16'hFFFF;
rommem[5594] <= 16'hFFFF;
rommem[5595] <= 16'hFFFF;
rommem[5596] <= 16'hFFFF;
rommem[5597] <= 16'hFFFF;
rommem[5598] <= 16'hFFFF;
rommem[5599] <= 16'hFFFF;
rommem[5600] <= 16'hFFFF;
rommem[5601] <= 16'hFFFF;
rommem[5602] <= 16'hFFFF;
rommem[5603] <= 16'hFFFF;
rommem[5604] <= 16'hFFFF;
rommem[5605] <= 16'hFFFF;
rommem[5606] <= 16'hFFFF;
rommem[5607] <= 16'hFFFF;
rommem[5608] <= 16'hFFFF;
rommem[5609] <= 16'hFFFF;
rommem[5610] <= 16'hFFFF;
rommem[5611] <= 16'hFFFF;
rommem[5612] <= 16'hFFFF;
rommem[5613] <= 16'hFFFF;
rommem[5614] <= 16'hFFFF;
rommem[5615] <= 16'hFFFF;
rommem[5616] <= 16'hFFFF;
rommem[5617] <= 16'hFFFF;
rommem[5618] <= 16'hFFFF;
rommem[5619] <= 16'hFFFF;
rommem[5620] <= 16'hFFFF;
rommem[5621] <= 16'hFFFF;
rommem[5622] <= 16'hFFFF;
rommem[5623] <= 16'hFFFF;
rommem[5624] <= 16'hFFFF;
rommem[5625] <= 16'hFFFF;
rommem[5626] <= 16'hFFFF;
rommem[5627] <= 16'hFFFF;
rommem[5628] <= 16'hFFFF;
rommem[5629] <= 16'hFFFF;
rommem[5630] <= 16'hFFFF;
rommem[5631] <= 16'hFFFF;
rommem[5632] <= 16'hFFFF;
rommem[5633] <= 16'hFFFF;
rommem[5634] <= 16'hFFFF;
rommem[5635] <= 16'hFFFF;
rommem[5636] <= 16'hFFFF;
rommem[5637] <= 16'hFFFF;
rommem[5638] <= 16'hFFFF;
rommem[5639] <= 16'hFFFF;
rommem[5640] <= 16'hFFFF;
rommem[5641] <= 16'hFFFF;
rommem[5642] <= 16'hFFFF;
rommem[5643] <= 16'hFFFF;
rommem[5644] <= 16'hFFFF;
rommem[5645] <= 16'hFFFF;
rommem[5646] <= 16'hFFFF;
rommem[5647] <= 16'hFFFF;
rommem[5648] <= 16'hFFFF;
rommem[5649] <= 16'hFFFF;
rommem[5650] <= 16'hFFFF;
rommem[5651] <= 16'hFFFF;
rommem[5652] <= 16'hFFFF;
rommem[5653] <= 16'hFFFF;
rommem[5654] <= 16'hFFFF;
rommem[5655] <= 16'hFFFF;
rommem[5656] <= 16'hFFFF;
rommem[5657] <= 16'hFFFF;
rommem[5658] <= 16'hFFFF;
rommem[5659] <= 16'hFFFF;
rommem[5660] <= 16'hFFFF;
rommem[5661] <= 16'hFFFF;
rommem[5662] <= 16'hFFFF;
rommem[5663] <= 16'hFFFF;
rommem[5664] <= 16'hFFFF;
rommem[5665] <= 16'hFFFF;
rommem[5666] <= 16'hFFFF;
rommem[5667] <= 16'hFFFF;
rommem[5668] <= 16'hFFFF;
rommem[5669] <= 16'hFFFF;
rommem[5670] <= 16'hFFFF;
rommem[5671] <= 16'hFFFF;
rommem[5672] <= 16'hFFFF;
rommem[5673] <= 16'hFFFF;
rommem[5674] <= 16'hFFFF;
rommem[5675] <= 16'hFFFF;
rommem[5676] <= 16'hFFFF;
rommem[5677] <= 16'hFFFF;
rommem[5678] <= 16'hFFFF;
rommem[5679] <= 16'hFFFF;
rommem[5680] <= 16'hFFFF;
rommem[5681] <= 16'hFFFF;
rommem[5682] <= 16'hFFFF;
rommem[5683] <= 16'hFFFF;
rommem[5684] <= 16'hFFFF;
rommem[5685] <= 16'hFFFF;
rommem[5686] <= 16'hFFFF;
rommem[5687] <= 16'hFFFF;
rommem[5688] <= 16'hFFFF;
rommem[5689] <= 16'hFFFF;
rommem[5690] <= 16'hFFFF;
rommem[5691] <= 16'hFFFF;
rommem[5692] <= 16'hFFFF;
rommem[5693] <= 16'hFFFF;
rommem[5694] <= 16'hFFFF;
rommem[5695] <= 16'hFFFF;
rommem[5696] <= 16'hFFFF;
rommem[5697] <= 16'hFFFF;
rommem[5698] <= 16'hFFFF;
rommem[5699] <= 16'hFFFF;
rommem[5700] <= 16'hFFFF;
rommem[5701] <= 16'hFFFF;
rommem[5702] <= 16'hFFFF;
rommem[5703] <= 16'hFFFF;
rommem[5704] <= 16'hFFFF;
rommem[5705] <= 16'hFFFF;
rommem[5706] <= 16'hFFFF;
rommem[5707] <= 16'hFFFF;
rommem[5708] <= 16'hFFFF;
rommem[5709] <= 16'hFFFF;
rommem[5710] <= 16'hFFFF;
rommem[5711] <= 16'hFFFF;
rommem[5712] <= 16'hFFFF;
rommem[5713] <= 16'hFFFF;
rommem[5714] <= 16'hFFFF;
rommem[5715] <= 16'hFFFF;
rommem[5716] <= 16'hFFFF;
rommem[5717] <= 16'hFFFF;
rommem[5718] <= 16'hFFFF;
rommem[5719] <= 16'hFFFF;
rommem[5720] <= 16'hFFFF;
rommem[5721] <= 16'hFFFF;
rommem[5722] <= 16'hFFFF;
rommem[5723] <= 16'hFFFF;
rommem[5724] <= 16'hFFFF;
rommem[5725] <= 16'hFFFF;
rommem[5726] <= 16'hFFFF;
rommem[5727] <= 16'hFFFF;
rommem[5728] <= 16'hFFFF;
rommem[5729] <= 16'hFFFF;
rommem[5730] <= 16'hFFFF;
rommem[5731] <= 16'hFFFF;
rommem[5732] <= 16'hFFFF;
rommem[5733] <= 16'hFFFF;
rommem[5734] <= 16'hFFFF;
rommem[5735] <= 16'hFFFF;
rommem[5736] <= 16'hFFFF;
rommem[5737] <= 16'hFFFF;
rommem[5738] <= 16'hFFFF;
rommem[5739] <= 16'hFFFF;
rommem[5740] <= 16'hFFFF;
rommem[5741] <= 16'hFFFF;
rommem[5742] <= 16'hFFFF;
rommem[5743] <= 16'hFFFF;
rommem[5744] <= 16'hFFFF;
rommem[5745] <= 16'hFFFF;
rommem[5746] <= 16'hFFFF;
rommem[5747] <= 16'hFFFF;
rommem[5748] <= 16'hFFFF;
rommem[5749] <= 16'hFFFF;
rommem[5750] <= 16'hFFFF;
rommem[5751] <= 16'hFFFF;
rommem[5752] <= 16'hFFFF;
rommem[5753] <= 16'hFFFF;
rommem[5754] <= 16'hFFFF;
rommem[5755] <= 16'hFFFF;
rommem[5756] <= 16'hFFFF;
rommem[5757] <= 16'hFFFF;
rommem[5758] <= 16'hFFFF;
rommem[5759] <= 16'hFFFF;
rommem[5760] <= 16'hFFFF;
rommem[5761] <= 16'hFFFF;
rommem[5762] <= 16'hFFFF;
rommem[5763] <= 16'hFFFF;
rommem[5764] <= 16'hFFFF;
rommem[5765] <= 16'hFFFF;
rommem[5766] <= 16'hFFFF;
rommem[5767] <= 16'hFFFF;
rommem[5768] <= 16'hFFFF;
rommem[5769] <= 16'hFFFF;
rommem[5770] <= 16'hFFFF;
rommem[5771] <= 16'hFFFF;
rommem[5772] <= 16'hFFFF;
rommem[5773] <= 16'hFFFF;
rommem[5774] <= 16'hFFFF;
rommem[5775] <= 16'hFFFF;
rommem[5776] <= 16'hFFFF;
rommem[5777] <= 16'hFFFF;
rommem[5778] <= 16'hFFFF;
rommem[5779] <= 16'hFFFF;
rommem[5780] <= 16'hFFFF;
rommem[5781] <= 16'hFFFF;
rommem[5782] <= 16'hFFFF;
rommem[5783] <= 16'hFFFF;
rommem[5784] <= 16'hFFFF;
rommem[5785] <= 16'hFFFF;
rommem[5786] <= 16'hFFFF;
rommem[5787] <= 16'hFFFF;
rommem[5788] <= 16'hFFFF;
rommem[5789] <= 16'hFFFF;
rommem[5790] <= 16'hFFFF;
rommem[5791] <= 16'hFFFF;
rommem[5792] <= 16'hFFFF;
rommem[5793] <= 16'hFFFF;
rommem[5794] <= 16'hFFFF;
rommem[5795] <= 16'hFFFF;
rommem[5796] <= 16'hFFFF;
rommem[5797] <= 16'hFFFF;
rommem[5798] <= 16'hFFFF;
rommem[5799] <= 16'hFFFF;
rommem[5800] <= 16'hFFFF;
rommem[5801] <= 16'hFFFF;
rommem[5802] <= 16'hFFFF;
rommem[5803] <= 16'hFFFF;
rommem[5804] <= 16'hFFFF;
rommem[5805] <= 16'hFFFF;
rommem[5806] <= 16'hFFFF;
rommem[5807] <= 16'hFFFF;
rommem[5808] <= 16'hFFFF;
rommem[5809] <= 16'hFFFF;
rommem[5810] <= 16'hFFFF;
rommem[5811] <= 16'hFFFF;
rommem[5812] <= 16'hFFFF;
rommem[5813] <= 16'hFFFF;
rommem[5814] <= 16'hFFFF;
rommem[5815] <= 16'hFFFF;
rommem[5816] <= 16'hFFFF;
rommem[5817] <= 16'hFFFF;
rommem[5818] <= 16'hFFFF;
rommem[5819] <= 16'hFFFF;
rommem[5820] <= 16'hFFFF;
rommem[5821] <= 16'hFFFF;
rommem[5822] <= 16'hFFFF;
rommem[5823] <= 16'hFFFF;
rommem[5824] <= 16'hFFFF;
rommem[5825] <= 16'hFFFF;
rommem[5826] <= 16'hFFFF;
rommem[5827] <= 16'hFFFF;
rommem[5828] <= 16'hFFFF;
rommem[5829] <= 16'hFFFF;
rommem[5830] <= 16'hFFFF;
rommem[5831] <= 16'hFFFF;
rommem[5832] <= 16'hFFFF;
rommem[5833] <= 16'hFFFF;
rommem[5834] <= 16'hFFFF;
rommem[5835] <= 16'hFFFF;
rommem[5836] <= 16'hFFFF;
rommem[5837] <= 16'hFFFF;
rommem[5838] <= 16'hFFFF;
rommem[5839] <= 16'hFFFF;
rommem[5840] <= 16'hFFFF;
rommem[5841] <= 16'hFFFF;
rommem[5842] <= 16'hFFFF;
rommem[5843] <= 16'hFFFF;
rommem[5844] <= 16'hFFFF;
rommem[5845] <= 16'hFFFF;
rommem[5846] <= 16'hFFFF;
rommem[5847] <= 16'hFFFF;
rommem[5848] <= 16'hFFFF;
rommem[5849] <= 16'hFFFF;
rommem[5850] <= 16'hFFFF;
rommem[5851] <= 16'hFFFF;
rommem[5852] <= 16'hFFFF;
rommem[5853] <= 16'hFFFF;
rommem[5854] <= 16'hFFFF;
rommem[5855] <= 16'hFFFF;
rommem[5856] <= 16'hFFFF;
rommem[5857] <= 16'hFFFF;
rommem[5858] <= 16'hFFFF;
rommem[5859] <= 16'hFFFF;
rommem[5860] <= 16'hFFFF;
rommem[5861] <= 16'hFFFF;
rommem[5862] <= 16'hFFFF;
rommem[5863] <= 16'hFFFF;
rommem[5864] <= 16'hFFFF;
rommem[5865] <= 16'hFFFF;
rommem[5866] <= 16'hFFFF;
rommem[5867] <= 16'hFFFF;
rommem[5868] <= 16'hFFFF;
rommem[5869] <= 16'hFFFF;
rommem[5870] <= 16'hFFFF;
rommem[5871] <= 16'hFFFF;
rommem[5872] <= 16'hFFFF;
rommem[5873] <= 16'hFFFF;
rommem[5874] <= 16'hFFFF;
rommem[5875] <= 16'hFFFF;
rommem[5876] <= 16'hFFFF;
rommem[5877] <= 16'hFFFF;
rommem[5878] <= 16'hFFFF;
rommem[5879] <= 16'hFFFF;
rommem[5880] <= 16'hFFFF;
rommem[5881] <= 16'hFFFF;
rommem[5882] <= 16'hFFFF;
rommem[5883] <= 16'hFFFF;
rommem[5884] <= 16'hFFFF;
rommem[5885] <= 16'hFFFF;
rommem[5886] <= 16'hFFFF;
rommem[5887] <= 16'hFFFF;
rommem[5888] <= 16'hFFFF;
rommem[5889] <= 16'hFFFF;
rommem[5890] <= 16'hFFFF;
rommem[5891] <= 16'hFFFF;
rommem[5892] <= 16'hFFFF;
rommem[5893] <= 16'hFFFF;
rommem[5894] <= 16'hFFFF;
rommem[5895] <= 16'hFFFF;
rommem[5896] <= 16'hFFFF;
rommem[5897] <= 16'hFFFF;
rommem[5898] <= 16'hFFFF;
rommem[5899] <= 16'hFFFF;
rommem[5900] <= 16'hFFFF;
rommem[5901] <= 16'hFFFF;
rommem[5902] <= 16'hFFFF;
rommem[5903] <= 16'hFFFF;
rommem[5904] <= 16'hFFFF;
rommem[5905] <= 16'hFFFF;
rommem[5906] <= 16'hFFFF;
rommem[5907] <= 16'hFFFF;
rommem[5908] <= 16'hFFFF;
rommem[5909] <= 16'hFFFF;
rommem[5910] <= 16'hFFFF;
rommem[5911] <= 16'hFFFF;
rommem[5912] <= 16'hFFFF;
rommem[5913] <= 16'hFFFF;
rommem[5914] <= 16'hFFFF;
rommem[5915] <= 16'hFFFF;
rommem[5916] <= 16'hFFFF;
rommem[5917] <= 16'hFFFF;
rommem[5918] <= 16'hFFFF;
rommem[5919] <= 16'hFFFF;
rommem[5920] <= 16'hFFFF;
rommem[5921] <= 16'hFFFF;
rommem[5922] <= 16'hFFFF;
rommem[5923] <= 16'hFFFF;
rommem[5924] <= 16'hFFFF;
rommem[5925] <= 16'hFFFF;
rommem[5926] <= 16'hFFFF;
rommem[5927] <= 16'hFFFF;
rommem[5928] <= 16'hFFFF;
rommem[5929] <= 16'hFFFF;
rommem[5930] <= 16'hFFFF;
rommem[5931] <= 16'hFFFF;
rommem[5932] <= 16'hFFFF;
rommem[5933] <= 16'hFFFF;
rommem[5934] <= 16'hFFFF;
rommem[5935] <= 16'hFFFF;
rommem[5936] <= 16'hFFFF;
rommem[5937] <= 16'hFFFF;
rommem[5938] <= 16'hFFFF;
rommem[5939] <= 16'hFFFF;
rommem[5940] <= 16'hFFFF;
rommem[5941] <= 16'hFFFF;
rommem[5942] <= 16'hFFFF;
rommem[5943] <= 16'hFFFF;
rommem[5944] <= 16'hFFFF;
rommem[5945] <= 16'hFFFF;
rommem[5946] <= 16'hFFFF;
rommem[5947] <= 16'hFFFF;
rommem[5948] <= 16'hFFFF;
rommem[5949] <= 16'hFFFF;
rommem[5950] <= 16'hFFFF;
rommem[5951] <= 16'hFFFF;
rommem[5952] <= 16'hFFFF;
rommem[5953] <= 16'hFFFF;
rommem[5954] <= 16'hFFFF;
rommem[5955] <= 16'hFFFF;
rommem[5956] <= 16'hFFFF;
rommem[5957] <= 16'hFFFF;
rommem[5958] <= 16'hFFFF;
rommem[5959] <= 16'hFFFF;
rommem[5960] <= 16'hFFFF;
rommem[5961] <= 16'hFFFF;
rommem[5962] <= 16'hFFFF;
rommem[5963] <= 16'hFFFF;
rommem[5964] <= 16'hFFFF;
rommem[5965] <= 16'hFFFF;
rommem[5966] <= 16'hFFFF;
rommem[5967] <= 16'hFFFF;
rommem[5968] <= 16'hFFFF;
rommem[5969] <= 16'hFFFF;
rommem[5970] <= 16'hFFFF;
rommem[5971] <= 16'hFFFF;
rommem[5972] <= 16'hFFFF;
rommem[5973] <= 16'hFFFF;
rommem[5974] <= 16'hFFFF;
rommem[5975] <= 16'hFFFF;
rommem[5976] <= 16'hFFFF;
rommem[5977] <= 16'hFFFF;
rommem[5978] <= 16'hFFFF;
rommem[5979] <= 16'hFFFF;
rommem[5980] <= 16'hFFFF;
rommem[5981] <= 16'hFFFF;
rommem[5982] <= 16'hFFFF;
rommem[5983] <= 16'hFFFF;
rommem[5984] <= 16'hFFFF;
rommem[5985] <= 16'hFFFF;
rommem[5986] <= 16'hFFFF;
rommem[5987] <= 16'hFFFF;
rommem[5988] <= 16'hFFFF;
rommem[5989] <= 16'hFFFF;
rommem[5990] <= 16'hFFFF;
rommem[5991] <= 16'hFFFF;
rommem[5992] <= 16'hFFFF;
rommem[5993] <= 16'hFFFF;
rommem[5994] <= 16'hFFFF;
rommem[5995] <= 16'hFFFF;
rommem[5996] <= 16'hFFFF;
rommem[5997] <= 16'hFFFF;
rommem[5998] <= 16'hFFFF;
rommem[5999] <= 16'hFFFF;
rommem[6000] <= 16'hFFFF;
rommem[6001] <= 16'hFFFF;
rommem[6002] <= 16'hFFFF;
rommem[6003] <= 16'hFFFF;
rommem[6004] <= 16'hFFFF;
rommem[6005] <= 16'hFFFF;
rommem[6006] <= 16'hFFFF;
rommem[6007] <= 16'hFFFF;
rommem[6008] <= 16'hFFFF;
rommem[6009] <= 16'hFFFF;
rommem[6010] <= 16'hFFFF;
rommem[6011] <= 16'hFFFF;
rommem[6012] <= 16'hFFFF;
rommem[6013] <= 16'hFFFF;
rommem[6014] <= 16'hFFFF;
rommem[6015] <= 16'hFFFF;
rommem[6016] <= 16'hFFFF;
rommem[6017] <= 16'hFFFF;
rommem[6018] <= 16'hFFFF;
rommem[6019] <= 16'hFFFF;
rommem[6020] <= 16'hFFFF;
rommem[6021] <= 16'hFFFF;
rommem[6022] <= 16'hFFFF;
rommem[6023] <= 16'hFFFF;
rommem[6024] <= 16'hFFFF;
rommem[6025] <= 16'hFFFF;
rommem[6026] <= 16'hFFFF;
rommem[6027] <= 16'hFFFF;
rommem[6028] <= 16'hFFFF;
rommem[6029] <= 16'hFFFF;
rommem[6030] <= 16'hFFFF;
rommem[6031] <= 16'hFFFF;
rommem[6032] <= 16'hFFFF;
rommem[6033] <= 16'hFFFF;
rommem[6034] <= 16'hFFFF;
rommem[6035] <= 16'hFFFF;
rommem[6036] <= 16'hFFFF;
rommem[6037] <= 16'hFFFF;
rommem[6038] <= 16'hFFFF;
rommem[6039] <= 16'hFFFF;
rommem[6040] <= 16'hFFFF;
rommem[6041] <= 16'hFFFF;
rommem[6042] <= 16'hFFFF;
rommem[6043] <= 16'hFFFF;
rommem[6044] <= 16'hFFFF;
rommem[6045] <= 16'hFFFF;
rommem[6046] <= 16'hFFFF;
rommem[6047] <= 16'hFFFF;
rommem[6048] <= 16'hFFFF;
rommem[6049] <= 16'hFFFF;
rommem[6050] <= 16'hFFFF;
rommem[6051] <= 16'hFFFF;
rommem[6052] <= 16'hFFFF;
rommem[6053] <= 16'hFFFF;
rommem[6054] <= 16'hFFFF;
rommem[6055] <= 16'hFFFF;
rommem[6056] <= 16'hFFFF;
rommem[6057] <= 16'hFFFF;
rommem[6058] <= 16'hFFFF;
rommem[6059] <= 16'hFFFF;
rommem[6060] <= 16'hFFFF;
rommem[6061] <= 16'hFFFF;
rommem[6062] <= 16'hFFFF;
rommem[6063] <= 16'hFFFF;
rommem[6064] <= 16'hFFFF;
rommem[6065] <= 16'hFFFF;
rommem[6066] <= 16'hFFFF;
rommem[6067] <= 16'hFFFF;
rommem[6068] <= 16'hFFFF;
rommem[6069] <= 16'hFFFF;
rommem[6070] <= 16'hFFFF;
rommem[6071] <= 16'hFFFF;
rommem[6072] <= 16'hFFFF;
rommem[6073] <= 16'hFFFF;
rommem[6074] <= 16'hFFFF;
rommem[6075] <= 16'hFFFF;
rommem[6076] <= 16'hFFFF;
rommem[6077] <= 16'hFFFF;
rommem[6078] <= 16'hFFFF;
rommem[6079] <= 16'hFFFF;
rommem[6080] <= 16'hFFFF;
rommem[6081] <= 16'hFFFF;
rommem[6082] <= 16'hFFFF;
rommem[6083] <= 16'hFFFF;
rommem[6084] <= 16'hFFFF;
rommem[6085] <= 16'hFFFF;
rommem[6086] <= 16'hFFFF;
rommem[6087] <= 16'hFFFF;
rommem[6088] <= 16'hFFFF;
rommem[6089] <= 16'hFFFF;
rommem[6090] <= 16'hFFFF;
rommem[6091] <= 16'hFFFF;
rommem[6092] <= 16'hFFFF;
rommem[6093] <= 16'hFFFF;
rommem[6094] <= 16'hFFFF;
rommem[6095] <= 16'hFFFF;
rommem[6096] <= 16'hFFFF;
rommem[6097] <= 16'hFFFF;
rommem[6098] <= 16'hFFFF;
rommem[6099] <= 16'hFFFF;
rommem[6100] <= 16'hFFFF;
rommem[6101] <= 16'hFFFF;
rommem[6102] <= 16'hFFFF;
rommem[6103] <= 16'hFFFF;
rommem[6104] <= 16'hFFFF;
rommem[6105] <= 16'hFFFF;
rommem[6106] <= 16'hFFFF;
rommem[6107] <= 16'hFFFF;
rommem[6108] <= 16'hFFFF;
rommem[6109] <= 16'hFFFF;
rommem[6110] <= 16'hFFFF;
rommem[6111] <= 16'hFFFF;
rommem[6112] <= 16'hFFFF;
rommem[6113] <= 16'hFFFF;
rommem[6114] <= 16'hFFFF;
rommem[6115] <= 16'hFFFF;
rommem[6116] <= 16'hFFFF;
rommem[6117] <= 16'hFFFF;
rommem[6118] <= 16'hFFFF;
rommem[6119] <= 16'hFFFF;
rommem[6120] <= 16'hFFFF;
rommem[6121] <= 16'hFFFF;
rommem[6122] <= 16'hFFFF;
rommem[6123] <= 16'hFFFF;
rommem[6124] <= 16'hFFFF;
rommem[6125] <= 16'hFFFF;
rommem[6126] <= 16'hFFFF;
rommem[6127] <= 16'hFFFF;
rommem[6128] <= 16'hFFFF;
rommem[6129] <= 16'hFFFF;
rommem[6130] <= 16'hFFFF;
rommem[6131] <= 16'hFFFF;
rommem[6132] <= 16'hFFFF;
rommem[6133] <= 16'hFFFF;
rommem[6134] <= 16'hFFFF;
rommem[6135] <= 16'hFFFF;
rommem[6136] <= 16'hFFFF;
rommem[6137] <= 16'hFFFF;
rommem[6138] <= 16'hFFFF;
rommem[6139] <= 16'hFFFF;
rommem[6140] <= 16'hFFFF;
rommem[6141] <= 16'hFFFF;
rommem[6142] <= 16'hFFFF;
rommem[6143] <= 16'hFFFF;
rommem[6144] <= 16'hFFFF;
rommem[6145] <= 16'hFFFF;
rommem[6146] <= 16'hFFFF;
rommem[6147] <= 16'hFFFF;
rommem[6148] <= 16'hFFFF;
rommem[6149] <= 16'hFFFF;
rommem[6150] <= 16'hFFFF;
rommem[6151] <= 16'hFFFF;
rommem[6152] <= 16'hFFFF;
rommem[6153] <= 16'hFFFF;
rommem[6154] <= 16'hFFFF;
rommem[6155] <= 16'hFFFF;
rommem[6156] <= 16'hFFFF;
rommem[6157] <= 16'hFFFF;
rommem[6158] <= 16'hFFFF;
rommem[6159] <= 16'hFFFF;
rommem[6160] <= 16'hFFFF;
rommem[6161] <= 16'hFFFF;
rommem[6162] <= 16'hFFFF;
rommem[6163] <= 16'hFFFF;
rommem[6164] <= 16'hFFFF;
rommem[6165] <= 16'hFFFF;
rommem[6166] <= 16'hFFFF;
rommem[6167] <= 16'hFFFF;
rommem[6168] <= 16'hFFFF;
rommem[6169] <= 16'hFFFF;
rommem[6170] <= 16'hFFFF;
rommem[6171] <= 16'hFFFF;
rommem[6172] <= 16'hFFFF;
rommem[6173] <= 16'hFFFF;
rommem[6174] <= 16'hFFFF;
rommem[6175] <= 16'hFFFF;
rommem[6176] <= 16'hFFFF;
rommem[6177] <= 16'hFFFF;
rommem[6178] <= 16'hFFFF;
rommem[6179] <= 16'hFFFF;
rommem[6180] <= 16'hFFFF;
rommem[6181] <= 16'hFFFF;
rommem[6182] <= 16'hFFFF;
rommem[6183] <= 16'hFFFF;
rommem[6184] <= 16'hFFFF;
rommem[6185] <= 16'hFFFF;
rommem[6186] <= 16'hFFFF;
rommem[6187] <= 16'hFFFF;
rommem[6188] <= 16'hFFFF;
rommem[6189] <= 16'hFFFF;
rommem[6190] <= 16'hFFFF;
rommem[6191] <= 16'hFFFF;
rommem[6192] <= 16'hFFFF;
rommem[6193] <= 16'hFFFF;
rommem[6194] <= 16'hFFFF;
rommem[6195] <= 16'hFFFF;
rommem[6196] <= 16'hFFFF;
rommem[6197] <= 16'hFFFF;
rommem[6198] <= 16'hFFFF;
rommem[6199] <= 16'hFFFF;
rommem[6200] <= 16'hFFFF;
rommem[6201] <= 16'hFFFF;
rommem[6202] <= 16'hFFFF;
rommem[6203] <= 16'hFFFF;
rommem[6204] <= 16'hFFFF;
rommem[6205] <= 16'hFFFF;
rommem[6206] <= 16'hFFFF;
rommem[6207] <= 16'hFFFF;
rommem[6208] <= 16'hFFFF;
rommem[6209] <= 16'hFFFF;
rommem[6210] <= 16'hFFFF;
rommem[6211] <= 16'hFFFF;
rommem[6212] <= 16'hFFFF;
rommem[6213] <= 16'hFFFF;
rommem[6214] <= 16'hFFFF;
rommem[6215] <= 16'hFFFF;
rommem[6216] <= 16'hFFFF;
rommem[6217] <= 16'hFFFF;
rommem[6218] <= 16'hFFFF;
rommem[6219] <= 16'hFFFF;
rommem[6220] <= 16'hFFFF;
rommem[6221] <= 16'hFFFF;
rommem[6222] <= 16'hFFFF;
rommem[6223] <= 16'hFFFF;
rommem[6224] <= 16'hFFFF;
rommem[6225] <= 16'hFFFF;
rommem[6226] <= 16'hFFFF;
rommem[6227] <= 16'hFFFF;
rommem[6228] <= 16'hFFFF;
rommem[6229] <= 16'hFFFF;
rommem[6230] <= 16'hFFFF;
rommem[6231] <= 16'hFFFF;
rommem[6232] <= 16'hFFFF;
rommem[6233] <= 16'hFFFF;
rommem[6234] <= 16'hFFFF;
rommem[6235] <= 16'hFFFF;
rommem[6236] <= 16'hFFFF;
rommem[6237] <= 16'hFFFF;
rommem[6238] <= 16'hFFFF;
rommem[6239] <= 16'hFFFF;
rommem[6240] <= 16'hFFFF;
rommem[6241] <= 16'hFFFF;
rommem[6242] <= 16'hFFFF;
rommem[6243] <= 16'hFFFF;
rommem[6244] <= 16'hFFFF;
rommem[6245] <= 16'hFFFF;
rommem[6246] <= 16'hFFFF;
rommem[6247] <= 16'hFFFF;
rommem[6248] <= 16'hFFFF;
rommem[6249] <= 16'hFFFF;
rommem[6250] <= 16'hFFFF;
rommem[6251] <= 16'hFFFF;
rommem[6252] <= 16'hFFFF;
rommem[6253] <= 16'hFFFF;
rommem[6254] <= 16'hFFFF;
rommem[6255] <= 16'hFFFF;
rommem[6256] <= 16'hFFFF;
rommem[6257] <= 16'hFFFF;
rommem[6258] <= 16'hFFFF;
rommem[6259] <= 16'hFFFF;
rommem[6260] <= 16'hFFFF;
rommem[6261] <= 16'hFFFF;
rommem[6262] <= 16'hFFFF;
rommem[6263] <= 16'hFFFF;
rommem[6264] <= 16'hFFFF;
rommem[6265] <= 16'hFFFF;
rommem[6266] <= 16'hFFFF;
rommem[6267] <= 16'hFFFF;
rommem[6268] <= 16'hFFFF;
rommem[6269] <= 16'hFFFF;
rommem[6270] <= 16'hFFFF;
rommem[6271] <= 16'hFFFF;
rommem[6272] <= 16'hFFFF;
rommem[6273] <= 16'hFFFF;
rommem[6274] <= 16'hFFFF;
rommem[6275] <= 16'hFFFF;
rommem[6276] <= 16'hFFFF;
rommem[6277] <= 16'hFFFF;
rommem[6278] <= 16'hFFFF;
rommem[6279] <= 16'hFFFF;
rommem[6280] <= 16'hFFFF;
rommem[6281] <= 16'hFFFF;
rommem[6282] <= 16'hFFFF;
rommem[6283] <= 16'hFFFF;
rommem[6284] <= 16'hFFFF;
rommem[6285] <= 16'hFFFF;
rommem[6286] <= 16'hFFFF;
rommem[6287] <= 16'hFFFF;
rommem[6288] <= 16'hFFFF;
rommem[6289] <= 16'hFFFF;
rommem[6290] <= 16'hFFFF;
rommem[6291] <= 16'hFFFF;
rommem[6292] <= 16'hFFFF;
rommem[6293] <= 16'hFFFF;
rommem[6294] <= 16'hFFFF;
rommem[6295] <= 16'hFFFF;
rommem[6296] <= 16'hFFFF;
rommem[6297] <= 16'hFFFF;
rommem[6298] <= 16'hFFFF;
rommem[6299] <= 16'hFFFF;
rommem[6300] <= 16'hFFFF;
rommem[6301] <= 16'hFFFF;
rommem[6302] <= 16'hFFFF;
rommem[6303] <= 16'hFFFF;
rommem[6304] <= 16'hFFFF;
rommem[6305] <= 16'hFFFF;
rommem[6306] <= 16'hFFFF;
rommem[6307] <= 16'hFFFF;
rommem[6308] <= 16'hFFFF;
rommem[6309] <= 16'hFFFF;
rommem[6310] <= 16'hFFFF;
rommem[6311] <= 16'hFFFF;
rommem[6312] <= 16'hFFFF;
rommem[6313] <= 16'hFFFF;
rommem[6314] <= 16'hFFFF;
rommem[6315] <= 16'hFFFF;
rommem[6316] <= 16'hFFFF;
rommem[6317] <= 16'hFFFF;
rommem[6318] <= 16'hFFFF;
rommem[6319] <= 16'hFFFF;
rommem[6320] <= 16'hFFFF;
rommem[6321] <= 16'hFFFF;
rommem[6322] <= 16'hFFFF;
rommem[6323] <= 16'hFFFF;
rommem[6324] <= 16'hFFFF;
rommem[6325] <= 16'hFFFF;
rommem[6326] <= 16'hFFFF;
rommem[6327] <= 16'hFFFF;
rommem[6328] <= 16'hFFFF;
rommem[6329] <= 16'hFFFF;
rommem[6330] <= 16'hFFFF;
rommem[6331] <= 16'hFFFF;
rommem[6332] <= 16'hFFFF;
rommem[6333] <= 16'hFFFF;
rommem[6334] <= 16'hFFFF;
rommem[6335] <= 16'hFFFF;
rommem[6336] <= 16'hFFFF;
rommem[6337] <= 16'hFFFF;
rommem[6338] <= 16'hFFFF;
rommem[6339] <= 16'hFFFF;
rommem[6340] <= 16'hFFFF;
rommem[6341] <= 16'hFFFF;
rommem[6342] <= 16'hFFFF;
rommem[6343] <= 16'hFFFF;
rommem[6344] <= 16'hFFFF;
rommem[6345] <= 16'hFFFF;
rommem[6346] <= 16'hFFFF;
rommem[6347] <= 16'hFFFF;
rommem[6348] <= 16'hFFFF;
rommem[6349] <= 16'hFFFF;
rommem[6350] <= 16'hFFFF;
rommem[6351] <= 16'hFFFF;
rommem[6352] <= 16'hFFFF;
rommem[6353] <= 16'hFFFF;
rommem[6354] <= 16'hFFFF;
rommem[6355] <= 16'hFFFF;
rommem[6356] <= 16'hFFFF;
rommem[6357] <= 16'hFFFF;
rommem[6358] <= 16'hFFFF;
rommem[6359] <= 16'hFFFF;
rommem[6360] <= 16'hFFFF;
rommem[6361] <= 16'hFFFF;
rommem[6362] <= 16'hFFFF;
rommem[6363] <= 16'hFFFF;
rommem[6364] <= 16'hFFFF;
rommem[6365] <= 16'hFFFF;
rommem[6366] <= 16'hFFFF;
rommem[6367] <= 16'hFFFF;
rommem[6368] <= 16'hFFFF;
rommem[6369] <= 16'hFFFF;
rommem[6370] <= 16'hFFFF;
rommem[6371] <= 16'hFFFF;
rommem[6372] <= 16'hFFFF;
rommem[6373] <= 16'hFFFF;
rommem[6374] <= 16'hFFFF;
rommem[6375] <= 16'hFFFF;
rommem[6376] <= 16'hFFFF;
rommem[6377] <= 16'hFFFF;
rommem[6378] <= 16'hFFFF;
rommem[6379] <= 16'hFFFF;
rommem[6380] <= 16'hFFFF;
rommem[6381] <= 16'hFFFF;
rommem[6382] <= 16'hFFFF;
rommem[6383] <= 16'hFFFF;
rommem[6384] <= 16'hFFFF;
rommem[6385] <= 16'hFFFF;
rommem[6386] <= 16'hFFFF;
rommem[6387] <= 16'hFFFF;
rommem[6388] <= 16'hFFFF;
rommem[6389] <= 16'hFFFF;
rommem[6390] <= 16'hFFFF;
rommem[6391] <= 16'hFFFF;
rommem[6392] <= 16'hFFFF;
rommem[6393] <= 16'hFFFF;
rommem[6394] <= 16'hFFFF;
rommem[6395] <= 16'hFFFF;
rommem[6396] <= 16'hFFFF;
rommem[6397] <= 16'hFFFF;
rommem[6398] <= 16'hFFFF;
rommem[6399] <= 16'hFFFF;
rommem[6400] <= 16'hFFFF;
rommem[6401] <= 16'hFFFF;
rommem[6402] <= 16'hFFFF;
rommem[6403] <= 16'hFFFF;
rommem[6404] <= 16'hFFFF;
rommem[6405] <= 16'hFFFF;
rommem[6406] <= 16'hFFFF;
rommem[6407] <= 16'hFFFF;
rommem[6408] <= 16'hFFFF;
rommem[6409] <= 16'hFFFF;
rommem[6410] <= 16'hFFFF;
rommem[6411] <= 16'hFFFF;
rommem[6412] <= 16'hFFFF;
rommem[6413] <= 16'hFFFF;
rommem[6414] <= 16'hFFFF;
rommem[6415] <= 16'hFFFF;
rommem[6416] <= 16'hFFFF;
rommem[6417] <= 16'hFFFF;
rommem[6418] <= 16'hFFFF;
rommem[6419] <= 16'hFFFF;
rommem[6420] <= 16'hFFFF;
rommem[6421] <= 16'hFFFF;
rommem[6422] <= 16'hFFFF;
rommem[6423] <= 16'hFFFF;
rommem[6424] <= 16'hFFFF;
rommem[6425] <= 16'hFFFF;
rommem[6426] <= 16'hFFFF;
rommem[6427] <= 16'hFFFF;
rommem[6428] <= 16'hFFFF;
rommem[6429] <= 16'hFFFF;
rommem[6430] <= 16'hFFFF;
rommem[6431] <= 16'hFFFF;
rommem[6432] <= 16'hFFFF;
rommem[6433] <= 16'hFFFF;
rommem[6434] <= 16'hFFFF;
rommem[6435] <= 16'hFFFF;
rommem[6436] <= 16'hFFFF;
rommem[6437] <= 16'hFFFF;
rommem[6438] <= 16'hFFFF;
rommem[6439] <= 16'hFFFF;
rommem[6440] <= 16'hFFFF;
rommem[6441] <= 16'hFFFF;
rommem[6442] <= 16'hFFFF;
rommem[6443] <= 16'hFFFF;
rommem[6444] <= 16'hFFFF;
rommem[6445] <= 16'hFFFF;
rommem[6446] <= 16'hFFFF;
rommem[6447] <= 16'hFFFF;
rommem[6448] <= 16'hFFFF;
rommem[6449] <= 16'hFFFF;
rommem[6450] <= 16'hFFFF;
rommem[6451] <= 16'hFFFF;
rommem[6452] <= 16'hFFFF;
rommem[6453] <= 16'hFFFF;
rommem[6454] <= 16'hFFFF;
rommem[6455] <= 16'hFFFF;
rommem[6456] <= 16'hFFFF;
rommem[6457] <= 16'hFFFF;
rommem[6458] <= 16'hFFFF;
rommem[6459] <= 16'hFFFF;
rommem[6460] <= 16'hFFFF;
rommem[6461] <= 16'hFFFF;
rommem[6462] <= 16'hFFFF;
rommem[6463] <= 16'hFFFF;
rommem[6464] <= 16'hFFFF;
rommem[6465] <= 16'hFFFF;
rommem[6466] <= 16'hFFFF;
rommem[6467] <= 16'hFFFF;
rommem[6468] <= 16'hFFFF;
rommem[6469] <= 16'hFFFF;
rommem[6470] <= 16'hFFFF;
rommem[6471] <= 16'hFFFF;
rommem[6472] <= 16'hFFFF;
rommem[6473] <= 16'hFFFF;
rommem[6474] <= 16'hFFFF;
rommem[6475] <= 16'hFFFF;
rommem[6476] <= 16'hFFFF;
rommem[6477] <= 16'hFFFF;
rommem[6478] <= 16'hFFFF;
rommem[6479] <= 16'hFFFF;
rommem[6480] <= 16'hFFFF;
rommem[6481] <= 16'hFFFF;
rommem[6482] <= 16'hFFFF;
rommem[6483] <= 16'hFFFF;
rommem[6484] <= 16'hFFFF;
rommem[6485] <= 16'hFFFF;
rommem[6486] <= 16'hFFFF;
rommem[6487] <= 16'hFFFF;
rommem[6488] <= 16'hFFFF;
rommem[6489] <= 16'hFFFF;
rommem[6490] <= 16'hFFFF;
rommem[6491] <= 16'hFFFF;
rommem[6492] <= 16'hFFFF;
rommem[6493] <= 16'hFFFF;
rommem[6494] <= 16'hFFFF;
rommem[6495] <= 16'hFFFF;
rommem[6496] <= 16'hFFFF;
rommem[6497] <= 16'hFFFF;
rommem[6498] <= 16'hFFFF;
rommem[6499] <= 16'hFFFF;
rommem[6500] <= 16'hFFFF;
rommem[6501] <= 16'hFFFF;
rommem[6502] <= 16'hFFFF;
rommem[6503] <= 16'hFFFF;
rommem[6504] <= 16'hFFFF;
rommem[6505] <= 16'hFFFF;
rommem[6506] <= 16'hFFFF;
rommem[6507] <= 16'hFFFF;
rommem[6508] <= 16'hFFFF;
rommem[6509] <= 16'hFFFF;
rommem[6510] <= 16'hFFFF;
rommem[6511] <= 16'hFFFF;
rommem[6512] <= 16'hFFFF;
rommem[6513] <= 16'hFFFF;
rommem[6514] <= 16'hFFFF;
rommem[6515] <= 16'hFFFF;
rommem[6516] <= 16'hFFFF;
rommem[6517] <= 16'hFFFF;
rommem[6518] <= 16'hFFFF;
rommem[6519] <= 16'hFFFF;
rommem[6520] <= 16'hFFFF;
rommem[6521] <= 16'hFFFF;
rommem[6522] <= 16'hFFFF;
rommem[6523] <= 16'hFFFF;
rommem[6524] <= 16'hFFFF;
rommem[6525] <= 16'hFFFF;
rommem[6526] <= 16'hFFFF;
rommem[6527] <= 16'hFFFF;
rommem[6528] <= 16'hFFFF;
rommem[6529] <= 16'hFFFF;
rommem[6530] <= 16'hFFFF;
rommem[6531] <= 16'hFFFF;
rommem[6532] <= 16'hFFFF;
rommem[6533] <= 16'hFFFF;
rommem[6534] <= 16'hFFFF;
rommem[6535] <= 16'hFFFF;
rommem[6536] <= 16'hFFFF;
rommem[6537] <= 16'hFFFF;
rommem[6538] <= 16'hFFFF;
rommem[6539] <= 16'hFFFF;
rommem[6540] <= 16'hFFFF;
rommem[6541] <= 16'hFFFF;
rommem[6542] <= 16'hFFFF;
rommem[6543] <= 16'hFFFF;
rommem[6544] <= 16'hFFFF;
rommem[6545] <= 16'hFFFF;
rommem[6546] <= 16'hFFFF;
rommem[6547] <= 16'hFFFF;
rommem[6548] <= 16'hFFFF;
rommem[6549] <= 16'hFFFF;
rommem[6550] <= 16'hFFFF;
rommem[6551] <= 16'hFFFF;
rommem[6552] <= 16'hFFFF;
rommem[6553] <= 16'hFFFF;
rommem[6554] <= 16'hFFFF;
rommem[6555] <= 16'hFFFF;
rommem[6556] <= 16'hFFFF;
rommem[6557] <= 16'hFFFF;
rommem[6558] <= 16'hFFFF;
rommem[6559] <= 16'hFFFF;
rommem[6560] <= 16'hFFFF;
rommem[6561] <= 16'hFFFF;
rommem[6562] <= 16'hFFFF;
rommem[6563] <= 16'hFFFF;
rommem[6564] <= 16'hFFFF;
rommem[6565] <= 16'hFFFF;
rommem[6566] <= 16'hFFFF;
rommem[6567] <= 16'hFFFF;
rommem[6568] <= 16'hFFFF;
rommem[6569] <= 16'hFFFF;
rommem[6570] <= 16'hFFFF;
rommem[6571] <= 16'hFFFF;
rommem[6572] <= 16'hFFFF;
rommem[6573] <= 16'hFFFF;
rommem[6574] <= 16'hFFFF;
rommem[6575] <= 16'hFFFF;
rommem[6576] <= 16'hFFFF;
rommem[6577] <= 16'hFFFF;
rommem[6578] <= 16'hFFFF;
rommem[6579] <= 16'hFFFF;
rommem[6580] <= 16'hFFFF;
rommem[6581] <= 16'hFFFF;
rommem[6582] <= 16'hFFFF;
rommem[6583] <= 16'hFFFF;
rommem[6584] <= 16'hFFFF;
rommem[6585] <= 16'hFFFF;
rommem[6586] <= 16'hFFFF;
rommem[6587] <= 16'hFFFF;
rommem[6588] <= 16'hFFFF;
rommem[6589] <= 16'hFFFF;
rommem[6590] <= 16'hFFFF;
rommem[6591] <= 16'hFFFF;
rommem[6592] <= 16'hFFFF;
rommem[6593] <= 16'hFFFF;
rommem[6594] <= 16'hFFFF;
rommem[6595] <= 16'hFFFF;
rommem[6596] <= 16'hFFFF;
rommem[6597] <= 16'hFFFF;
rommem[6598] <= 16'hFFFF;
rommem[6599] <= 16'hFFFF;
rommem[6600] <= 16'hFFFF;
rommem[6601] <= 16'hFFFF;
rommem[6602] <= 16'hFFFF;
rommem[6603] <= 16'hFFFF;
rommem[6604] <= 16'hFFFF;
rommem[6605] <= 16'hFFFF;
rommem[6606] <= 16'hFFFF;
rommem[6607] <= 16'hFFFF;
rommem[6608] <= 16'hFFFF;
rommem[6609] <= 16'hFFFF;
rommem[6610] <= 16'hFFFF;
rommem[6611] <= 16'hFFFF;
rommem[6612] <= 16'hFFFF;
rommem[6613] <= 16'hFFFF;
rommem[6614] <= 16'hFFFF;
rommem[6615] <= 16'hFFFF;
rommem[6616] <= 16'hFFFF;
rommem[6617] <= 16'hFFFF;
rommem[6618] <= 16'hFFFF;
rommem[6619] <= 16'hFFFF;
rommem[6620] <= 16'hFFFF;
rommem[6621] <= 16'hFFFF;
rommem[6622] <= 16'hFFFF;
rommem[6623] <= 16'hFFFF;
rommem[6624] <= 16'hFFFF;
rommem[6625] <= 16'hFFFF;
rommem[6626] <= 16'hFFFF;
rommem[6627] <= 16'hFFFF;
rommem[6628] <= 16'hFFFF;
rommem[6629] <= 16'hFFFF;
rommem[6630] <= 16'hFFFF;
rommem[6631] <= 16'hFFFF;
rommem[6632] <= 16'hFFFF;
rommem[6633] <= 16'hFFFF;
rommem[6634] <= 16'hFFFF;
rommem[6635] <= 16'hFFFF;
rommem[6636] <= 16'hFFFF;
rommem[6637] <= 16'hFFFF;
rommem[6638] <= 16'hFFFF;
rommem[6639] <= 16'hFFFF;
rommem[6640] <= 16'hFFFF;
rommem[6641] <= 16'hFFFF;
rommem[6642] <= 16'hFFFF;
rommem[6643] <= 16'hFFFF;
rommem[6644] <= 16'hFFFF;
rommem[6645] <= 16'hFFFF;
rommem[6646] <= 16'hFFFF;
rommem[6647] <= 16'hFFFF;
rommem[6648] <= 16'hFFFF;
rommem[6649] <= 16'hFFFF;
rommem[6650] <= 16'hFFFF;
rommem[6651] <= 16'hFFFF;
rommem[6652] <= 16'hFFFF;
rommem[6653] <= 16'hFFFF;
rommem[6654] <= 16'hFFFF;
rommem[6655] <= 16'hFFFF;
rommem[6656] <= 16'hFFFF;
rommem[6657] <= 16'hFFFF;
rommem[6658] <= 16'hFFFF;
rommem[6659] <= 16'hFFFF;
rommem[6660] <= 16'hFFFF;
rommem[6661] <= 16'hFFFF;
rommem[6662] <= 16'hFFFF;
rommem[6663] <= 16'hFFFF;
rommem[6664] <= 16'hFFFF;
rommem[6665] <= 16'hFFFF;
rommem[6666] <= 16'hFFFF;
rommem[6667] <= 16'hFFFF;
rommem[6668] <= 16'hFFFF;
rommem[6669] <= 16'hFFFF;
rommem[6670] <= 16'hFFFF;
rommem[6671] <= 16'hFFFF;
rommem[6672] <= 16'hFFFF;
rommem[6673] <= 16'hFFFF;
rommem[6674] <= 16'hFFFF;
rommem[6675] <= 16'hFFFF;
rommem[6676] <= 16'hFFFF;
rommem[6677] <= 16'hFFFF;
rommem[6678] <= 16'hFFFF;
rommem[6679] <= 16'hFFFF;
rommem[6680] <= 16'hFFFF;
rommem[6681] <= 16'hFFFF;
rommem[6682] <= 16'hFFFF;
rommem[6683] <= 16'hFFFF;
rommem[6684] <= 16'hFFFF;
rommem[6685] <= 16'hFFFF;
rommem[6686] <= 16'hFFFF;
rommem[6687] <= 16'hFFFF;
rommem[6688] <= 16'hFFFF;
rommem[6689] <= 16'hFFFF;
rommem[6690] <= 16'hFFFF;
rommem[6691] <= 16'hFFFF;
rommem[6692] <= 16'hFFFF;
rommem[6693] <= 16'hFFFF;
rommem[6694] <= 16'hFFFF;
rommem[6695] <= 16'hFFFF;
rommem[6696] <= 16'hFFFF;
rommem[6697] <= 16'hFFFF;
rommem[6698] <= 16'hFFFF;
rommem[6699] <= 16'hFFFF;
rommem[6700] <= 16'hFFFF;
rommem[6701] <= 16'hFFFF;
rommem[6702] <= 16'hFFFF;
rommem[6703] <= 16'hFFFF;
rommem[6704] <= 16'hFFFF;
rommem[6705] <= 16'hFFFF;
rommem[6706] <= 16'hFFFF;
rommem[6707] <= 16'hFFFF;
rommem[6708] <= 16'hFFFF;
rommem[6709] <= 16'hFFFF;
rommem[6710] <= 16'hFFFF;
rommem[6711] <= 16'hFFFF;
rommem[6712] <= 16'hFFFF;
rommem[6713] <= 16'hFFFF;
rommem[6714] <= 16'hFFFF;
rommem[6715] <= 16'hFFFF;
rommem[6716] <= 16'hFFFF;
rommem[6717] <= 16'hFFFF;
rommem[6718] <= 16'hFFFF;
rommem[6719] <= 16'hFFFF;
rommem[6720] <= 16'hFFFF;
rommem[6721] <= 16'hFFFF;
rommem[6722] <= 16'hFFFF;
rommem[6723] <= 16'hFFFF;
rommem[6724] <= 16'hFFFF;
rommem[6725] <= 16'hFFFF;
rommem[6726] <= 16'hFFFF;
rommem[6727] <= 16'hFFFF;
rommem[6728] <= 16'hFFFF;
rommem[6729] <= 16'hFFFF;
rommem[6730] <= 16'hFFFF;
rommem[6731] <= 16'hFFFF;
rommem[6732] <= 16'hFFFF;
rommem[6733] <= 16'hFFFF;
rommem[6734] <= 16'hFFFF;
rommem[6735] <= 16'hFFFF;
rommem[6736] <= 16'hFFFF;
rommem[6737] <= 16'hFFFF;
rommem[6738] <= 16'hFFFF;
rommem[6739] <= 16'hFFFF;
rommem[6740] <= 16'hFFFF;
rommem[6741] <= 16'hFFFF;
rommem[6742] <= 16'hFFFF;
rommem[6743] <= 16'hFFFF;
rommem[6744] <= 16'hFFFF;
rommem[6745] <= 16'hFFFF;
rommem[6746] <= 16'hFFFF;
rommem[6747] <= 16'hFFFF;
rommem[6748] <= 16'hFFFF;
rommem[6749] <= 16'hFFFF;
rommem[6750] <= 16'hFFFF;
rommem[6751] <= 16'hFFFF;
rommem[6752] <= 16'hFFFF;
rommem[6753] <= 16'hFFFF;
rommem[6754] <= 16'hFFFF;
rommem[6755] <= 16'hFFFF;
rommem[6756] <= 16'hFFFF;
rommem[6757] <= 16'hFFFF;
rommem[6758] <= 16'hFFFF;
rommem[6759] <= 16'hFFFF;
rommem[6760] <= 16'hFFFF;
rommem[6761] <= 16'hFFFF;
rommem[6762] <= 16'hFFFF;
rommem[6763] <= 16'hFFFF;
rommem[6764] <= 16'hFFFF;
rommem[6765] <= 16'hFFFF;
rommem[6766] <= 16'hFFFF;
rommem[6767] <= 16'hFFFF;
rommem[6768] <= 16'hFFFF;
rommem[6769] <= 16'hFFFF;
rommem[6770] <= 16'hFFFF;
rommem[6771] <= 16'hFFFF;
rommem[6772] <= 16'hFFFF;
rommem[6773] <= 16'hFFFF;
rommem[6774] <= 16'hFFFF;
rommem[6775] <= 16'hFFFF;
rommem[6776] <= 16'hFFFF;
rommem[6777] <= 16'hFFFF;
rommem[6778] <= 16'hFFFF;
rommem[6779] <= 16'hFFFF;
rommem[6780] <= 16'hFFFF;
rommem[6781] <= 16'hFFFF;
rommem[6782] <= 16'hFFFF;
rommem[6783] <= 16'hFFFF;
rommem[6784] <= 16'hFFFF;
rommem[6785] <= 16'hFFFF;
rommem[6786] <= 16'hFFFF;
rommem[6787] <= 16'hFFFF;
rommem[6788] <= 16'hFFFF;
rommem[6789] <= 16'hFFFF;
rommem[6790] <= 16'hFFFF;
rommem[6791] <= 16'hFFFF;
rommem[6792] <= 16'hFFFF;
rommem[6793] <= 16'hFFFF;
rommem[6794] <= 16'hFFFF;
rommem[6795] <= 16'hFFFF;
rommem[6796] <= 16'hFFFF;
rommem[6797] <= 16'hFFFF;
rommem[6798] <= 16'hFFFF;
rommem[6799] <= 16'hFFFF;
rommem[6800] <= 16'hFFFF;
rommem[6801] <= 16'hFFFF;
rommem[6802] <= 16'hFFFF;
rommem[6803] <= 16'hFFFF;
rommem[6804] <= 16'hFFFF;
rommem[6805] <= 16'hFFFF;
rommem[6806] <= 16'hFFFF;
rommem[6807] <= 16'hFFFF;
rommem[6808] <= 16'hFFFF;
rommem[6809] <= 16'hFFFF;
rommem[6810] <= 16'hFFFF;
rommem[6811] <= 16'hFFFF;
rommem[6812] <= 16'hFFFF;
rommem[6813] <= 16'hFFFF;
rommem[6814] <= 16'hFFFF;
rommem[6815] <= 16'hFFFF;
rommem[6816] <= 16'hFFFF;
rommem[6817] <= 16'hFFFF;
rommem[6818] <= 16'hFFFF;
rommem[6819] <= 16'hFFFF;
rommem[6820] <= 16'hFFFF;
rommem[6821] <= 16'hFFFF;
rommem[6822] <= 16'hFFFF;
rommem[6823] <= 16'hFFFF;
rommem[6824] <= 16'hFFFF;
rommem[6825] <= 16'hFFFF;
rommem[6826] <= 16'hFFFF;
rommem[6827] <= 16'hFFFF;
rommem[6828] <= 16'hFFFF;
rommem[6829] <= 16'hFFFF;
rommem[6830] <= 16'hFFFF;
rommem[6831] <= 16'hFFFF;
rommem[6832] <= 16'hFFFF;
rommem[6833] <= 16'hFFFF;
rommem[6834] <= 16'hFFFF;
rommem[6835] <= 16'hFFFF;
rommem[6836] <= 16'hFFFF;
rommem[6837] <= 16'hFFFF;
rommem[6838] <= 16'hFFFF;
rommem[6839] <= 16'hFFFF;
rommem[6840] <= 16'hFFFF;
rommem[6841] <= 16'hFFFF;
rommem[6842] <= 16'hFFFF;
rommem[6843] <= 16'hFFFF;
rommem[6844] <= 16'hFFFF;
rommem[6845] <= 16'hFFFF;
rommem[6846] <= 16'hFFFF;
rommem[6847] <= 16'hFFFF;
rommem[6848] <= 16'hFFFF;
rommem[6849] <= 16'hFFFF;
rommem[6850] <= 16'hFFFF;
rommem[6851] <= 16'hFFFF;
rommem[6852] <= 16'hFFFF;
rommem[6853] <= 16'hFFFF;
rommem[6854] <= 16'hFFFF;
rommem[6855] <= 16'hFFFF;
rommem[6856] <= 16'hFFFF;
rommem[6857] <= 16'hFFFF;
rommem[6858] <= 16'hFFFF;
rommem[6859] <= 16'hFFFF;
rommem[6860] <= 16'hFFFF;
rommem[6861] <= 16'hFFFF;
rommem[6862] <= 16'hFFFF;
rommem[6863] <= 16'hFFFF;
rommem[6864] <= 16'hFFFF;
rommem[6865] <= 16'hFFFF;
rommem[6866] <= 16'hFFFF;
rommem[6867] <= 16'hFFFF;
rommem[6868] <= 16'hFFFF;
rommem[6869] <= 16'hFFFF;
rommem[6870] <= 16'hFFFF;
rommem[6871] <= 16'hFFFF;
rommem[6872] <= 16'hFFFF;
rommem[6873] <= 16'hFFFF;
rommem[6874] <= 16'hFFFF;
rommem[6875] <= 16'hFFFF;
rommem[6876] <= 16'hFFFF;
rommem[6877] <= 16'hFFFF;
rommem[6878] <= 16'hFFFF;
rommem[6879] <= 16'hFFFF;
rommem[6880] <= 16'hFFFF;
rommem[6881] <= 16'hFFFF;
rommem[6882] <= 16'hFFFF;
rommem[6883] <= 16'hFFFF;
rommem[6884] <= 16'hFFFF;
rommem[6885] <= 16'hFFFF;
rommem[6886] <= 16'hFFFF;
rommem[6887] <= 16'hFFFF;
rommem[6888] <= 16'hFFFF;
rommem[6889] <= 16'hFFFF;
rommem[6890] <= 16'hFFFF;
rommem[6891] <= 16'hFFFF;
rommem[6892] <= 16'hFFFF;
rommem[6893] <= 16'hFFFF;
rommem[6894] <= 16'hFFFF;
rommem[6895] <= 16'hFFFF;
rommem[6896] <= 16'hFFFF;
rommem[6897] <= 16'hFFFF;
rommem[6898] <= 16'hFFFF;
rommem[6899] <= 16'hFFFF;
rommem[6900] <= 16'hFFFF;
rommem[6901] <= 16'hFFFF;
rommem[6902] <= 16'hFFFF;
rommem[6903] <= 16'hFFFF;
rommem[6904] <= 16'hFFFF;
rommem[6905] <= 16'hFFFF;
rommem[6906] <= 16'hFFFF;
rommem[6907] <= 16'hFFFF;
rommem[6908] <= 16'hFFFF;
rommem[6909] <= 16'hFFFF;
rommem[6910] <= 16'hFFFF;
rommem[6911] <= 16'hFFFF;
rommem[6912] <= 16'hFFFF;
rommem[6913] <= 16'hFFFF;
rommem[6914] <= 16'hFFFF;
rommem[6915] <= 16'hFFFF;
rommem[6916] <= 16'hFFFF;
rommem[6917] <= 16'hFFFF;
rommem[6918] <= 16'hFFFF;
rommem[6919] <= 16'hFFFF;
rommem[6920] <= 16'hFFFF;
rommem[6921] <= 16'hFFFF;
rommem[6922] <= 16'hFFFF;
rommem[6923] <= 16'hFFFF;
rommem[6924] <= 16'hFFFF;
rommem[6925] <= 16'hFFFF;
rommem[6926] <= 16'hFFFF;
rommem[6927] <= 16'hFFFF;
rommem[6928] <= 16'hFFFF;
rommem[6929] <= 16'hFFFF;
rommem[6930] <= 16'hFFFF;
rommem[6931] <= 16'hFFFF;
rommem[6932] <= 16'hFFFF;
rommem[6933] <= 16'hFFFF;
rommem[6934] <= 16'hFFFF;
rommem[6935] <= 16'hFFFF;
rommem[6936] <= 16'hFFFF;
rommem[6937] <= 16'hFFFF;
rommem[6938] <= 16'hFFFF;
rommem[6939] <= 16'hFFFF;
rommem[6940] <= 16'hFFFF;
rommem[6941] <= 16'hFFFF;
rommem[6942] <= 16'hFFFF;
rommem[6943] <= 16'hFFFF;
rommem[6944] <= 16'hFFFF;
rommem[6945] <= 16'hFFFF;
rommem[6946] <= 16'hFFFF;
rommem[6947] <= 16'hFFFF;
rommem[6948] <= 16'hFFFF;
rommem[6949] <= 16'hFFFF;
rommem[6950] <= 16'hFFFF;
rommem[6951] <= 16'hFFFF;
rommem[6952] <= 16'hFFFF;
rommem[6953] <= 16'hFFFF;
rommem[6954] <= 16'hFFFF;
rommem[6955] <= 16'hFFFF;
rommem[6956] <= 16'hFFFF;
rommem[6957] <= 16'hFFFF;
rommem[6958] <= 16'hFFFF;
rommem[6959] <= 16'hFFFF;
rommem[6960] <= 16'hFFFF;
rommem[6961] <= 16'hFFFF;
rommem[6962] <= 16'hFFFF;
rommem[6963] <= 16'hFFFF;
rommem[6964] <= 16'hFFFF;
rommem[6965] <= 16'hFFFF;
rommem[6966] <= 16'hFFFF;
rommem[6967] <= 16'hFFFF;
rommem[6968] <= 16'hFFFF;
rommem[6969] <= 16'hFFFF;
rommem[6970] <= 16'hFFFF;
rommem[6971] <= 16'hFFFF;
rommem[6972] <= 16'hFFFF;
rommem[6973] <= 16'hFFFF;
rommem[6974] <= 16'hFFFF;
rommem[6975] <= 16'hFFFF;
rommem[6976] <= 16'hFFFF;
rommem[6977] <= 16'hFFFF;
rommem[6978] <= 16'hFFFF;
rommem[6979] <= 16'hFFFF;
rommem[6980] <= 16'hFFFF;
rommem[6981] <= 16'hFFFF;
rommem[6982] <= 16'hFFFF;
rommem[6983] <= 16'hFFFF;
rommem[6984] <= 16'hFFFF;
rommem[6985] <= 16'hFFFF;
rommem[6986] <= 16'hFFFF;
rommem[6987] <= 16'hFFFF;
rommem[6988] <= 16'hFFFF;
rommem[6989] <= 16'hFFFF;
rommem[6990] <= 16'hFFFF;
rommem[6991] <= 16'hFFFF;
rommem[6992] <= 16'hFFFF;
rommem[6993] <= 16'hFFFF;
rommem[6994] <= 16'hFFFF;
rommem[6995] <= 16'hFFFF;
rommem[6996] <= 16'hFFFF;
rommem[6997] <= 16'hFFFF;
rommem[6998] <= 16'hFFFF;
rommem[6999] <= 16'hFFFF;
rommem[7000] <= 16'hFFFF;
rommem[7001] <= 16'hFFFF;
rommem[7002] <= 16'hFFFF;
rommem[7003] <= 16'hFFFF;
rommem[7004] <= 16'hFFFF;
rommem[7005] <= 16'hFFFF;
rommem[7006] <= 16'hFFFF;
rommem[7007] <= 16'hFFFF;
rommem[7008] <= 16'hFFFF;
rommem[7009] <= 16'hFFFF;
rommem[7010] <= 16'hFFFF;
rommem[7011] <= 16'hFFFF;
rommem[7012] <= 16'hFFFF;
rommem[7013] <= 16'hFFFF;
rommem[7014] <= 16'hFFFF;
rommem[7015] <= 16'hFFFF;
rommem[7016] <= 16'hFFFF;
rommem[7017] <= 16'hFFFF;
rommem[7018] <= 16'hFFFF;
rommem[7019] <= 16'hFFFF;
rommem[7020] <= 16'hFFFF;
rommem[7021] <= 16'hFFFF;
rommem[7022] <= 16'hFFFF;
rommem[7023] <= 16'hFFFF;
rommem[7024] <= 16'hFFFF;
rommem[7025] <= 16'hFFFF;
rommem[7026] <= 16'hFFFF;
rommem[7027] <= 16'hFFFF;
rommem[7028] <= 16'hFFFF;
rommem[7029] <= 16'hFFFF;
rommem[7030] <= 16'hFFFF;
rommem[7031] <= 16'hFFFF;
rommem[7032] <= 16'hFFFF;
rommem[7033] <= 16'hFFFF;
rommem[7034] <= 16'hFFFF;
rommem[7035] <= 16'hFFFF;
rommem[7036] <= 16'hFFFF;
rommem[7037] <= 16'hFFFF;
rommem[7038] <= 16'hFFFF;
rommem[7039] <= 16'hFFFF;
rommem[7040] <= 16'hFFFF;
rommem[7041] <= 16'hFFFF;
rommem[7042] <= 16'hFFFF;
rommem[7043] <= 16'hFFFF;
rommem[7044] <= 16'hFFFF;
rommem[7045] <= 16'hFFFF;
rommem[7046] <= 16'hFFFF;
rommem[7047] <= 16'hFFFF;
rommem[7048] <= 16'hFFFF;
rommem[7049] <= 16'hFFFF;
rommem[7050] <= 16'hFFFF;
rommem[7051] <= 16'hFFFF;
rommem[7052] <= 16'hFFFF;
rommem[7053] <= 16'hFFFF;
rommem[7054] <= 16'hFFFF;
rommem[7055] <= 16'hFFFF;
rommem[7056] <= 16'hFFFF;
rommem[7057] <= 16'hFFFF;
rommem[7058] <= 16'hFFFF;
rommem[7059] <= 16'hFFFF;
rommem[7060] <= 16'hFFFF;
rommem[7061] <= 16'hFFFF;
rommem[7062] <= 16'hFFFF;
rommem[7063] <= 16'hFFFF;
rommem[7064] <= 16'hFFFF;
rommem[7065] <= 16'hFFFF;
rommem[7066] <= 16'hFFFF;
rommem[7067] <= 16'hFFFF;
rommem[7068] <= 16'hFFFF;
rommem[7069] <= 16'hFFFF;
rommem[7070] <= 16'hFFFF;
rommem[7071] <= 16'hFFFF;
rommem[7072] <= 16'hFFFF;
rommem[7073] <= 16'hFFFF;
rommem[7074] <= 16'hFFFF;
rommem[7075] <= 16'hFFFF;
rommem[7076] <= 16'hFFFF;
rommem[7077] <= 16'hFFFF;
rommem[7078] <= 16'hFFFF;
rommem[7079] <= 16'hFFFF;
rommem[7080] <= 16'hFFFF;
rommem[7081] <= 16'hFFFF;
rommem[7082] <= 16'hFFFF;
rommem[7083] <= 16'hFFFF;
rommem[7084] <= 16'hFFFF;
rommem[7085] <= 16'hFFFF;
rommem[7086] <= 16'hFFFF;
rommem[7087] <= 16'hFFFF;
rommem[7088] <= 16'hFFFF;
rommem[7089] <= 16'hFFFF;
rommem[7090] <= 16'hFFFF;
rommem[7091] <= 16'hFFFF;
rommem[7092] <= 16'hFFFF;
rommem[7093] <= 16'hFFFF;
rommem[7094] <= 16'hFFFF;
rommem[7095] <= 16'hFFFF;
rommem[7096] <= 16'hFFFF;
rommem[7097] <= 16'hFFFF;
rommem[7098] <= 16'hFFFF;
rommem[7099] <= 16'hFFFF;
rommem[7100] <= 16'hFFFF;
rommem[7101] <= 16'hFFFF;
rommem[7102] <= 16'hFFFF;
rommem[7103] <= 16'hFFFF;
rommem[7104] <= 16'hFFFF;
rommem[7105] <= 16'hFFFF;
rommem[7106] <= 16'hFFFF;
rommem[7107] <= 16'hFFFF;
rommem[7108] <= 16'hFFFF;
rommem[7109] <= 16'hFFFF;
rommem[7110] <= 16'hFFFF;
rommem[7111] <= 16'hFFFF;
rommem[7112] <= 16'hFFFF;
rommem[7113] <= 16'hFFFF;
rommem[7114] <= 16'hFFFF;
rommem[7115] <= 16'hFFFF;
rommem[7116] <= 16'hFFFF;
rommem[7117] <= 16'hFFFF;
rommem[7118] <= 16'hFFFF;
rommem[7119] <= 16'hFFFF;
rommem[7120] <= 16'hFFFF;
rommem[7121] <= 16'hFFFF;
rommem[7122] <= 16'hFFFF;
rommem[7123] <= 16'hFFFF;
rommem[7124] <= 16'hFFFF;
rommem[7125] <= 16'hFFFF;
rommem[7126] <= 16'hFFFF;
rommem[7127] <= 16'hFFFF;
rommem[7128] <= 16'hFFFF;
rommem[7129] <= 16'hFFFF;
rommem[7130] <= 16'hFFFF;
rommem[7131] <= 16'hFFFF;
rommem[7132] <= 16'hFFFF;
rommem[7133] <= 16'hFFFF;
rommem[7134] <= 16'hFFFF;
rommem[7135] <= 16'hFFFF;
rommem[7136] <= 16'hFFFF;
rommem[7137] <= 16'hFFFF;
rommem[7138] <= 16'hFFFF;
rommem[7139] <= 16'hFFFF;
rommem[7140] <= 16'hFFFF;
rommem[7141] <= 16'hFFFF;
rommem[7142] <= 16'hFFFF;
rommem[7143] <= 16'hFFFF;
rommem[7144] <= 16'hFFFF;
rommem[7145] <= 16'hFFFF;
rommem[7146] <= 16'hFFFF;
rommem[7147] <= 16'hFFFF;
rommem[7148] <= 16'hFFFF;
rommem[7149] <= 16'hFFFF;
rommem[7150] <= 16'hFFFF;
rommem[7151] <= 16'hFFFF;
rommem[7152] <= 16'hFFFF;
rommem[7153] <= 16'hFFFF;
rommem[7154] <= 16'hFFFF;
rommem[7155] <= 16'hFFFF;
rommem[7156] <= 16'hFFFF;
rommem[7157] <= 16'hFFFF;
rommem[7158] <= 16'hFFFF;
rommem[7159] <= 16'hFFFF;
rommem[7160] <= 16'hFFFF;
rommem[7161] <= 16'hFFFF;
rommem[7162] <= 16'hFFFF;
rommem[7163] <= 16'hFFFF;
rommem[7164] <= 16'hFFFF;
rommem[7165] <= 16'hFFFF;
rommem[7166] <= 16'hFFFF;
rommem[7167] <= 16'hFFFF;
rommem[7168] <= 16'hFFFF;
rommem[7169] <= 16'hFFFF;
rommem[7170] <= 16'hFFFF;
rommem[7171] <= 16'hFFFF;
rommem[7172] <= 16'hFFFF;
rommem[7173] <= 16'hFFFF;
rommem[7174] <= 16'hFFFF;
rommem[7175] <= 16'hFFFF;
rommem[7176] <= 16'hFFFF;
rommem[7177] <= 16'hFFFF;
rommem[7178] <= 16'hFFFF;
rommem[7179] <= 16'hFFFF;
rommem[7180] <= 16'hFFFF;
rommem[7181] <= 16'hFFFF;
rommem[7182] <= 16'hFFFF;
rommem[7183] <= 16'hFFFF;
rommem[7184] <= 16'hFFFF;
rommem[7185] <= 16'hFFFF;
rommem[7186] <= 16'hFFFF;
rommem[7187] <= 16'hFFFF;
rommem[7188] <= 16'hFFFF;
rommem[7189] <= 16'hFFFF;
rommem[7190] <= 16'hFFFF;
rommem[7191] <= 16'hFFFF;
rommem[7192] <= 16'hFFFF;
rommem[7193] <= 16'hFFFF;
rommem[7194] <= 16'hFFFF;
rommem[7195] <= 16'hFFFF;
rommem[7196] <= 16'hFFFF;
rommem[7197] <= 16'hFFFF;
rommem[7198] <= 16'hFFFF;
rommem[7199] <= 16'hFFFF;
rommem[7200] <= 16'hFFFF;
rommem[7201] <= 16'hFFFF;
rommem[7202] <= 16'hFFFF;
rommem[7203] <= 16'hFFFF;
rommem[7204] <= 16'hFFFF;
rommem[7205] <= 16'hFFFF;
rommem[7206] <= 16'hFFFF;
rommem[7207] <= 16'hFFFF;
rommem[7208] <= 16'hFFFF;
rommem[7209] <= 16'hFFFF;
rommem[7210] <= 16'hFFFF;
rommem[7211] <= 16'hFFFF;
rommem[7212] <= 16'hFFFF;
rommem[7213] <= 16'hFFFF;
rommem[7214] <= 16'hFFFF;
rommem[7215] <= 16'hFFFF;
rommem[7216] <= 16'hFFFF;
rommem[7217] <= 16'hFFFF;
rommem[7218] <= 16'hFFFF;
rommem[7219] <= 16'hFFFF;
rommem[7220] <= 16'hFFFF;
rommem[7221] <= 16'hFFFF;
rommem[7222] <= 16'hFFFF;
rommem[7223] <= 16'hFFFF;
rommem[7224] <= 16'hFFFF;
rommem[7225] <= 16'hFFFF;
rommem[7226] <= 16'hFFFF;
rommem[7227] <= 16'hFFFF;
rommem[7228] <= 16'hFFFF;
rommem[7229] <= 16'hFFFF;
rommem[7230] <= 16'hFFFF;
rommem[7231] <= 16'hFFFF;
rommem[7232] <= 16'hFFFF;
rommem[7233] <= 16'hFFFF;
rommem[7234] <= 16'hFFFF;
rommem[7235] <= 16'hFFFF;
rommem[7236] <= 16'hFFFF;
rommem[7237] <= 16'hFFFF;
rommem[7238] <= 16'hFFFF;
rommem[7239] <= 16'hFFFF;
rommem[7240] <= 16'hFFFF;
rommem[7241] <= 16'hFFFF;
rommem[7242] <= 16'hFFFF;
rommem[7243] <= 16'hFFFF;
rommem[7244] <= 16'hFFFF;
rommem[7245] <= 16'hFFFF;
rommem[7246] <= 16'hFFFF;
rommem[7247] <= 16'hFFFF;
rommem[7248] <= 16'hFFFF;
rommem[7249] <= 16'hFFFF;
rommem[7250] <= 16'hFFFF;
rommem[7251] <= 16'hFFFF;
rommem[7252] <= 16'hFFFF;
rommem[7253] <= 16'hFFFF;
rommem[7254] <= 16'hFFFF;
rommem[7255] <= 16'hFFFF;
rommem[7256] <= 16'hFFFF;
rommem[7257] <= 16'hFFFF;
rommem[7258] <= 16'hFFFF;
rommem[7259] <= 16'hFFFF;
rommem[7260] <= 16'hFFFF;
rommem[7261] <= 16'hFFFF;
rommem[7262] <= 16'hFFFF;
rommem[7263] <= 16'hFFFF;
rommem[7264] <= 16'hFFFF;
rommem[7265] <= 16'hFFFF;
rommem[7266] <= 16'hFFFF;
rommem[7267] <= 16'hFFFF;
rommem[7268] <= 16'hFFFF;
rommem[7269] <= 16'hFFFF;
rommem[7270] <= 16'hFFFF;
rommem[7271] <= 16'hFFFF;
rommem[7272] <= 16'hFFFF;
rommem[7273] <= 16'hFFFF;
rommem[7274] <= 16'hFFFF;
rommem[7275] <= 16'hFFFF;
rommem[7276] <= 16'hFFFF;
rommem[7277] <= 16'hFFFF;
rommem[7278] <= 16'hFFFF;
rommem[7279] <= 16'hFFFF;
rommem[7280] <= 16'hFFFF;
rommem[7281] <= 16'hFFFF;
rommem[7282] <= 16'hFFFF;
rommem[7283] <= 16'hFFFF;
rommem[7284] <= 16'hFFFF;
rommem[7285] <= 16'hFFFF;
rommem[7286] <= 16'hFFFF;
rommem[7287] <= 16'hFFFF;
rommem[7288] <= 16'hFFFF;
rommem[7289] <= 16'hFFFF;
rommem[7290] <= 16'hFFFF;
rommem[7291] <= 16'hFFFF;
rommem[7292] <= 16'hFFFF;
rommem[7293] <= 16'hFFFF;
rommem[7294] <= 16'hFFFF;
rommem[7295] <= 16'hFFFF;
rommem[7296] <= 16'hFFFF;
rommem[7297] <= 16'hFFFF;
rommem[7298] <= 16'hFFFF;
rommem[7299] <= 16'hFFFF;
rommem[7300] <= 16'hFFFF;
rommem[7301] <= 16'hFFFF;
rommem[7302] <= 16'hFFFF;
rommem[7303] <= 16'hFFFF;
rommem[7304] <= 16'hFFFF;
rommem[7305] <= 16'hFFFF;
rommem[7306] <= 16'hFFFF;
rommem[7307] <= 16'hFFFF;
rommem[7308] <= 16'hFFFF;
rommem[7309] <= 16'hFFFF;
rommem[7310] <= 16'hFFFF;
rommem[7311] <= 16'hFFFF;
rommem[7312] <= 16'hFFFF;
rommem[7313] <= 16'hFFFF;
rommem[7314] <= 16'hFFFF;
rommem[7315] <= 16'hFFFF;
rommem[7316] <= 16'hFFFF;
rommem[7317] <= 16'hFFFF;
rommem[7318] <= 16'hFFFF;
rommem[7319] <= 16'hFFFF;
rommem[7320] <= 16'hFFFF;
rommem[7321] <= 16'hFFFF;
rommem[7322] <= 16'hFFFF;
rommem[7323] <= 16'hFFFF;
rommem[7324] <= 16'hFFFF;
rommem[7325] <= 16'hFFFF;
rommem[7326] <= 16'hFFFF;
rommem[7327] <= 16'hFFFF;
rommem[7328] <= 16'hFFFF;
rommem[7329] <= 16'hFFFF;
rommem[7330] <= 16'hFFFF;
rommem[7331] <= 16'hFFFF;
rommem[7332] <= 16'hFFFF;
rommem[7333] <= 16'hFFFF;
rommem[7334] <= 16'hFFFF;
rommem[7335] <= 16'hFFFF;
rommem[7336] <= 16'hFFFF;
rommem[7337] <= 16'hFFFF;
rommem[7338] <= 16'hFFFF;
rommem[7339] <= 16'hFFFF;
rommem[7340] <= 16'hFFFF;
rommem[7341] <= 16'hFFFF;
rommem[7342] <= 16'hFFFF;
rommem[7343] <= 16'hFFFF;
rommem[7344] <= 16'hFFFF;
rommem[7345] <= 16'hFFFF;
rommem[7346] <= 16'hFFFF;
rommem[7347] <= 16'hFFFF;
rommem[7348] <= 16'hFFFF;
rommem[7349] <= 16'hFFFF;
rommem[7350] <= 16'hFFFF;
rommem[7351] <= 16'hFFFF;
rommem[7352] <= 16'hFFFF;
rommem[7353] <= 16'hFFFF;
rommem[7354] <= 16'hFFFF;
rommem[7355] <= 16'hFFFF;
rommem[7356] <= 16'hFFFF;
rommem[7357] <= 16'hFFFF;
rommem[7358] <= 16'hFFFF;
rommem[7359] <= 16'hFFFF;
rommem[7360] <= 16'hFFFF;
rommem[7361] <= 16'hFFFF;
rommem[7362] <= 16'hFFFF;
rommem[7363] <= 16'hFFFF;
rommem[7364] <= 16'hFFFF;
rommem[7365] <= 16'hFFFF;
rommem[7366] <= 16'hFFFF;
rommem[7367] <= 16'hFFFF;
rommem[7368] <= 16'hFFFF;
rommem[7369] <= 16'hFFFF;
rommem[7370] <= 16'hFFFF;
rommem[7371] <= 16'hFFFF;
rommem[7372] <= 16'hFFFF;
rommem[7373] <= 16'hFFFF;
rommem[7374] <= 16'hFFFF;
rommem[7375] <= 16'hFFFF;
rommem[7376] <= 16'hFFFF;
rommem[7377] <= 16'hFFFF;
rommem[7378] <= 16'hFFFF;
rommem[7379] <= 16'hFFFF;
rommem[7380] <= 16'hFFFF;
rommem[7381] <= 16'hFFFF;
rommem[7382] <= 16'hFFFF;
rommem[7383] <= 16'hFFFF;
rommem[7384] <= 16'hFFFF;
rommem[7385] <= 16'hFFFF;
rommem[7386] <= 16'hFFFF;
rommem[7387] <= 16'hFFFF;
rommem[7388] <= 16'hFFFF;
rommem[7389] <= 16'hFFFF;
rommem[7390] <= 16'hFFFF;
rommem[7391] <= 16'hFFFF;
rommem[7392] <= 16'hFFFF;
rommem[7393] <= 16'hFFFF;
rommem[7394] <= 16'hFFFF;
rommem[7395] <= 16'hFFFF;
rommem[7396] <= 16'hFFFF;
rommem[7397] <= 16'hFFFF;
rommem[7398] <= 16'hFFFF;
rommem[7399] <= 16'hFFFF;
rommem[7400] <= 16'hFFFF;
rommem[7401] <= 16'hFFFF;
rommem[7402] <= 16'hFFFF;
rommem[7403] <= 16'hFFFF;
rommem[7404] <= 16'hFFFF;
rommem[7405] <= 16'hFFFF;
rommem[7406] <= 16'hFFFF;
rommem[7407] <= 16'hFFFF;
rommem[7408] <= 16'hFFFF;
rommem[7409] <= 16'hFFFF;
rommem[7410] <= 16'hFFFF;
rommem[7411] <= 16'hFFFF;
rommem[7412] <= 16'hFFFF;
rommem[7413] <= 16'hFFFF;
rommem[7414] <= 16'hFFFF;
rommem[7415] <= 16'hFFFF;
rommem[7416] <= 16'hFFFF;
rommem[7417] <= 16'hFFFF;
rommem[7418] <= 16'hFFFF;
rommem[7419] <= 16'hFFFF;
rommem[7420] <= 16'hFFFF;
rommem[7421] <= 16'hFFFF;
rommem[7422] <= 16'hFFFF;
rommem[7423] <= 16'hFFFF;
rommem[7424] <= 16'hFFFF;
rommem[7425] <= 16'hFFFF;
rommem[7426] <= 16'hFFFF;
rommem[7427] <= 16'hFFFF;
rommem[7428] <= 16'hFFFF;
rommem[7429] <= 16'hFFFF;
rommem[7430] <= 16'hFFFF;
rommem[7431] <= 16'hFFFF;
rommem[7432] <= 16'hFFFF;
rommem[7433] <= 16'hFFFF;
rommem[7434] <= 16'hFFFF;
rommem[7435] <= 16'hFFFF;
rommem[7436] <= 16'hFFFF;
rommem[7437] <= 16'hFFFF;
rommem[7438] <= 16'hFFFF;
rommem[7439] <= 16'hFFFF;
rommem[7440] <= 16'hFFFF;
rommem[7441] <= 16'hFFFF;
rommem[7442] <= 16'hFFFF;
rommem[7443] <= 16'hFFFF;
rommem[7444] <= 16'hFFFF;
rommem[7445] <= 16'hFFFF;
rommem[7446] <= 16'hFFFF;
rommem[7447] <= 16'hFFFF;
rommem[7448] <= 16'hFFFF;
rommem[7449] <= 16'hFFFF;
rommem[7450] <= 16'hFFFF;
rommem[7451] <= 16'hFFFF;
rommem[7452] <= 16'hFFFF;
rommem[7453] <= 16'hFFFF;
rommem[7454] <= 16'hFFFF;
rommem[7455] <= 16'hFFFF;
rommem[7456] <= 16'hFFFF;
rommem[7457] <= 16'hFFFF;
rommem[7458] <= 16'hFFFF;
rommem[7459] <= 16'hFFFF;
rommem[7460] <= 16'hFFFF;
rommem[7461] <= 16'hFFFF;
rommem[7462] <= 16'hFFFF;
rommem[7463] <= 16'hFFFF;
rommem[7464] <= 16'hFFFF;
rommem[7465] <= 16'hFFFF;
rommem[7466] <= 16'hFFFF;
rommem[7467] <= 16'hFFFF;
rommem[7468] <= 16'hFFFF;
rommem[7469] <= 16'hFFFF;
rommem[7470] <= 16'hFFFF;
rommem[7471] <= 16'hFFFF;
rommem[7472] <= 16'hFFFF;
rommem[7473] <= 16'hFFFF;
rommem[7474] <= 16'hFFFF;
rommem[7475] <= 16'hFFFF;
rommem[7476] <= 16'hFFFF;
rommem[7477] <= 16'hFFFF;
rommem[7478] <= 16'hFFFF;
rommem[7479] <= 16'hFFFF;
rommem[7480] <= 16'hFFFF;
rommem[7481] <= 16'hFFFF;
rommem[7482] <= 16'hFFFF;
rommem[7483] <= 16'hFFFF;
rommem[7484] <= 16'hFFFF;
rommem[7485] <= 16'hFFFF;
rommem[7486] <= 16'hFFFF;
rommem[7487] <= 16'hFFFF;
rommem[7488] <= 16'hFFFF;
rommem[7489] <= 16'hFFFF;
rommem[7490] <= 16'hFFFF;
rommem[7491] <= 16'hFFFF;
rommem[7492] <= 16'hFFFF;
rommem[7493] <= 16'hFFFF;
rommem[7494] <= 16'hFFFF;
rommem[7495] <= 16'hFFFF;
rommem[7496] <= 16'hFFFF;
rommem[7497] <= 16'hFFFF;
rommem[7498] <= 16'hFFFF;
rommem[7499] <= 16'hFFFF;
rommem[7500] <= 16'hFFFF;
rommem[7501] <= 16'hFFFF;
rommem[7502] <= 16'hFFFF;
rommem[7503] <= 16'hFFFF;
rommem[7504] <= 16'hFFFF;
rommem[7505] <= 16'hFFFF;
rommem[7506] <= 16'hFFFF;
rommem[7507] <= 16'hFFFF;
rommem[7508] <= 16'hFFFF;
rommem[7509] <= 16'hFFFF;
rommem[7510] <= 16'hFFFF;
rommem[7511] <= 16'hFFFF;
rommem[7512] <= 16'hFFFF;
rommem[7513] <= 16'hFFFF;
rommem[7514] <= 16'hFFFF;
rommem[7515] <= 16'hFFFF;
rommem[7516] <= 16'hFFFF;
rommem[7517] <= 16'hFFFF;
rommem[7518] <= 16'hFFFF;
rommem[7519] <= 16'hFFFF;
rommem[7520] <= 16'hFFFF;
rommem[7521] <= 16'hFFFF;
rommem[7522] <= 16'hFFFF;
rommem[7523] <= 16'hFFFF;
rommem[7524] <= 16'hFFFF;
rommem[7525] <= 16'hFFFF;
rommem[7526] <= 16'hFFFF;
rommem[7527] <= 16'hFFFF;
rommem[7528] <= 16'hFFFF;
rommem[7529] <= 16'hFFFF;
rommem[7530] <= 16'hFFFF;
rommem[7531] <= 16'hFFFF;
rommem[7532] <= 16'hFFFF;
rommem[7533] <= 16'hFFFF;
rommem[7534] <= 16'hFFFF;
rommem[7535] <= 16'hFFFF;
rommem[7536] <= 16'hFFFF;
rommem[7537] <= 16'hFFFF;
rommem[7538] <= 16'hFFFF;
rommem[7539] <= 16'hFFFF;
rommem[7540] <= 16'hFFFF;
rommem[7541] <= 16'hFFFF;
rommem[7542] <= 16'hFFFF;
rommem[7543] <= 16'hFFFF;
rommem[7544] <= 16'hFFFF;
rommem[7545] <= 16'hFFFF;
rommem[7546] <= 16'hFFFF;
rommem[7547] <= 16'hFFFF;
rommem[7548] <= 16'hFFFF;
rommem[7549] <= 16'hFFFF;
rommem[7550] <= 16'hFFFF;
rommem[7551] <= 16'hFFFF;
rommem[7552] <= 16'hFFFF;
rommem[7553] <= 16'hFFFF;
rommem[7554] <= 16'hFFFF;
rommem[7555] <= 16'hFFFF;
rommem[7556] <= 16'hFFFF;
rommem[7557] <= 16'hFFFF;
rommem[7558] <= 16'hFFFF;
rommem[7559] <= 16'hFFFF;
rommem[7560] <= 16'hFFFF;
rommem[7561] <= 16'hFFFF;
rommem[7562] <= 16'hFFFF;
rommem[7563] <= 16'hFFFF;
rommem[7564] <= 16'hFFFF;
rommem[7565] <= 16'hFFFF;
rommem[7566] <= 16'hFFFF;
rommem[7567] <= 16'hFFFF;
rommem[7568] <= 16'hFFFF;
rommem[7569] <= 16'hFFFF;
rommem[7570] <= 16'hFFFF;
rommem[7571] <= 16'hFFFF;
rommem[7572] <= 16'hFFFF;
rommem[7573] <= 16'hFFFF;
rommem[7574] <= 16'hFFFF;
rommem[7575] <= 16'hFFFF;
rommem[7576] <= 16'hFFFF;
rommem[7577] <= 16'hFFFF;
rommem[7578] <= 16'hFFFF;
rommem[7579] <= 16'hFFFF;
rommem[7580] <= 16'hFFFF;
rommem[7581] <= 16'hFFFF;
rommem[7582] <= 16'hFFFF;
rommem[7583] <= 16'hFFFF;
rommem[7584] <= 16'hFFFF;
rommem[7585] <= 16'hFFFF;
rommem[7586] <= 16'hFFFF;
rommem[7587] <= 16'hFFFF;
rommem[7588] <= 16'hFFFF;
rommem[7589] <= 16'hFFFF;
rommem[7590] <= 16'hFFFF;
rommem[7591] <= 16'hFFFF;
rommem[7592] <= 16'hFFFF;
rommem[7593] <= 16'hFFFF;
rommem[7594] <= 16'hFFFF;
rommem[7595] <= 16'hFFFF;
rommem[7596] <= 16'hFFFF;
rommem[7597] <= 16'hFFFF;
rommem[7598] <= 16'hFFFF;
rommem[7599] <= 16'hFFFF;
rommem[7600] <= 16'hFFFF;
rommem[7601] <= 16'hFFFF;
rommem[7602] <= 16'hFFFF;
rommem[7603] <= 16'hFFFF;
rommem[7604] <= 16'hFFFF;
rommem[7605] <= 16'hFFFF;
rommem[7606] <= 16'hFFFF;
rommem[7607] <= 16'hFFFF;
rommem[7608] <= 16'hFFFF;
rommem[7609] <= 16'hFFFF;
rommem[7610] <= 16'hFFFF;
rommem[7611] <= 16'hFFFF;
rommem[7612] <= 16'hFFFF;
rommem[7613] <= 16'hFFFF;
rommem[7614] <= 16'hFFFF;
rommem[7615] <= 16'hFFFF;
rommem[7616] <= 16'hFFFF;
rommem[7617] <= 16'hFFFF;
rommem[7618] <= 16'hFFFF;
rommem[7619] <= 16'hFFFF;
rommem[7620] <= 16'hFFFF;
rommem[7621] <= 16'hFFFF;
rommem[7622] <= 16'hFFFF;
rommem[7623] <= 16'hFFFF;
rommem[7624] <= 16'hFFFF;
rommem[7625] <= 16'hFFFF;
rommem[7626] <= 16'hFFFF;
rommem[7627] <= 16'hFFFF;
rommem[7628] <= 16'hFFFF;
rommem[7629] <= 16'hFFFF;
rommem[7630] <= 16'hFFFF;
rommem[7631] <= 16'hFFFF;
rommem[7632] <= 16'hFFFF;
rommem[7633] <= 16'hFFFF;
rommem[7634] <= 16'hFFFF;
rommem[7635] <= 16'hFFFF;
rommem[7636] <= 16'hFFFF;
rommem[7637] <= 16'hFFFF;
rommem[7638] <= 16'hFFFF;
rommem[7639] <= 16'hFFFF;
rommem[7640] <= 16'hFFFF;
rommem[7641] <= 16'hFFFF;
rommem[7642] <= 16'hFFFF;
rommem[7643] <= 16'hFFFF;
rommem[7644] <= 16'hFFFF;
rommem[7645] <= 16'hFFFF;
rommem[7646] <= 16'hFFFF;
rommem[7647] <= 16'hFFFF;
rommem[7648] <= 16'hFFFF;
rommem[7649] <= 16'hFFFF;
rommem[7650] <= 16'hFFFF;
rommem[7651] <= 16'hFFFF;
rommem[7652] <= 16'hFFFF;
rommem[7653] <= 16'hFFFF;
rommem[7654] <= 16'hFFFF;
rommem[7655] <= 16'hFFFF;
rommem[7656] <= 16'hFFFF;
rommem[7657] <= 16'hFFFF;
rommem[7658] <= 16'hFFFF;
rommem[7659] <= 16'hFFFF;
rommem[7660] <= 16'hFFFF;
rommem[7661] <= 16'hFFFF;
rommem[7662] <= 16'hFFFF;
rommem[7663] <= 16'hFFFF;
rommem[7664] <= 16'hFFFF;
rommem[7665] <= 16'hFFFF;
rommem[7666] <= 16'hFFFF;
rommem[7667] <= 16'hFFFF;
rommem[7668] <= 16'hFFFF;
rommem[7669] <= 16'hFFFF;
rommem[7670] <= 16'hFFFF;
rommem[7671] <= 16'hFFFF;
rommem[7672] <= 16'hFFFF;
rommem[7673] <= 16'hFFFF;
rommem[7674] <= 16'hFFFF;
rommem[7675] <= 16'hFFFF;
rommem[7676] <= 16'hFFFF;
rommem[7677] <= 16'hFFFF;
rommem[7678] <= 16'hFFFF;
rommem[7679] <= 16'hFFFF;
rommem[7680] <= 16'hFFFF;
rommem[7681] <= 16'hFFFF;
rommem[7682] <= 16'hFFFF;
rommem[7683] <= 16'hFFFF;
rommem[7684] <= 16'hFFFF;
rommem[7685] <= 16'hFFFF;
rommem[7686] <= 16'hFFFF;
rommem[7687] <= 16'hFFFF;
rommem[7688] <= 16'hFFFF;
rommem[7689] <= 16'hFFFF;
rommem[7690] <= 16'hFFFF;
rommem[7691] <= 16'hFFFF;
rommem[7692] <= 16'hFFFF;
rommem[7693] <= 16'hFFFF;
rommem[7694] <= 16'hFFFF;
rommem[7695] <= 16'hFFFF;
rommem[7696] <= 16'hFFFF;
rommem[7697] <= 16'hFFFF;
rommem[7698] <= 16'hFFFF;
rommem[7699] <= 16'hFFFF;
rommem[7700] <= 16'hFFFF;
rommem[7701] <= 16'hFFFF;
rommem[7702] <= 16'hFFFF;
rommem[7703] <= 16'hFFFF;
rommem[7704] <= 16'hFFFF;
rommem[7705] <= 16'hFFFF;
rommem[7706] <= 16'hFFFF;
rommem[7707] <= 16'hFFFF;
rommem[7708] <= 16'hFFFF;
rommem[7709] <= 16'hFFFF;
rommem[7710] <= 16'hFFFF;
rommem[7711] <= 16'hFFFF;
rommem[7712] <= 16'hFFFF;
rommem[7713] <= 16'hFFFF;
rommem[7714] <= 16'hFFFF;
rommem[7715] <= 16'hFFFF;
rommem[7716] <= 16'hFFFF;
rommem[7717] <= 16'hFFFF;
rommem[7718] <= 16'hFFFF;
rommem[7719] <= 16'hFFFF;
rommem[7720] <= 16'hFFFF;
rommem[7721] <= 16'hFFFF;
rommem[7722] <= 16'hFFFF;
rommem[7723] <= 16'hFFFF;
rommem[7724] <= 16'hFFFF;
rommem[7725] <= 16'hFFFF;
rommem[7726] <= 16'hFFFF;
rommem[7727] <= 16'hFFFF;
rommem[7728] <= 16'hFFFF;
rommem[7729] <= 16'hFFFF;
rommem[7730] <= 16'hFFFF;
rommem[7731] <= 16'hFFFF;
rommem[7732] <= 16'hFFFF;
rommem[7733] <= 16'hFFFF;
rommem[7734] <= 16'hFFFF;
rommem[7735] <= 16'hFFFF;
rommem[7736] <= 16'hFFFF;
rommem[7737] <= 16'hFFFF;
rommem[7738] <= 16'hFFFF;
rommem[7739] <= 16'hFFFF;
rommem[7740] <= 16'hFFFF;
rommem[7741] <= 16'hFFFF;
rommem[7742] <= 16'hFFFF;
rommem[7743] <= 16'hFFFF;
rommem[7744] <= 16'hFFFF;
rommem[7745] <= 16'hFFFF;
rommem[7746] <= 16'hFFFF;
rommem[7747] <= 16'hFFFF;
rommem[7748] <= 16'hFFFF;
rommem[7749] <= 16'hFFFF;
rommem[7750] <= 16'hFFFF;
rommem[7751] <= 16'hFFFF;
rommem[7752] <= 16'hFFFF;
rommem[7753] <= 16'hFFFF;
rommem[7754] <= 16'hFFFF;
rommem[7755] <= 16'hFFFF;
rommem[7756] <= 16'hFFFF;
rommem[7757] <= 16'hFFFF;
rommem[7758] <= 16'hFFFF;
rommem[7759] <= 16'hFFFF;
rommem[7760] <= 16'hFFFF;
rommem[7761] <= 16'hFFFF;
rommem[7762] <= 16'hFFFF;
rommem[7763] <= 16'hFFFF;
rommem[7764] <= 16'hFFFF;
rommem[7765] <= 16'hFFFF;
rommem[7766] <= 16'hFFFF;
rommem[7767] <= 16'hFFFF;
rommem[7768] <= 16'hFFFF;
rommem[7769] <= 16'hFFFF;
rommem[7770] <= 16'hFFFF;
rommem[7771] <= 16'hFFFF;
rommem[7772] <= 16'hFFFF;
rommem[7773] <= 16'hFFFF;
rommem[7774] <= 16'hFFFF;
rommem[7775] <= 16'hFFFF;
rommem[7776] <= 16'hFFFF;
rommem[7777] <= 16'hFFFF;
rommem[7778] <= 16'hFFFF;
rommem[7779] <= 16'hFFFF;
rommem[7780] <= 16'hFFFF;
rommem[7781] <= 16'hFFFF;
rommem[7782] <= 16'hFFFF;
rommem[7783] <= 16'hFFFF;
rommem[7784] <= 16'hFFFF;
rommem[7785] <= 16'hFFFF;
rommem[7786] <= 16'hFFFF;
rommem[7787] <= 16'hFFFF;
rommem[7788] <= 16'hFFFF;
rommem[7789] <= 16'hFFFF;
rommem[7790] <= 16'hFFFF;
rommem[7791] <= 16'hFFFF;
rommem[7792] <= 16'hFFFF;
rommem[7793] <= 16'hFFFF;
rommem[7794] <= 16'hFFFF;
rommem[7795] <= 16'hFFFF;
rommem[7796] <= 16'hFFFF;
rommem[7797] <= 16'hFFFF;
rommem[7798] <= 16'hFFFF;
rommem[7799] <= 16'hFFFF;
rommem[7800] <= 16'hFFFF;
rommem[7801] <= 16'hFFFF;
rommem[7802] <= 16'hFFFF;
rommem[7803] <= 16'hFFFF;
rommem[7804] <= 16'hFFFF;
rommem[7805] <= 16'hFFFF;
rommem[7806] <= 16'hFFFF;
rommem[7807] <= 16'hFFFF;
rommem[7808] <= 16'hFFFF;
rommem[7809] <= 16'hFFFF;
rommem[7810] <= 16'hFFFF;
rommem[7811] <= 16'hFFFF;
rommem[7812] <= 16'hFFFF;
rommem[7813] <= 16'hFFFF;
rommem[7814] <= 16'hFFFF;
rommem[7815] <= 16'hFFFF;
rommem[7816] <= 16'hFFFF;
rommem[7817] <= 16'hFFFF;
rommem[7818] <= 16'hFFFF;
rommem[7819] <= 16'hFFFF;
rommem[7820] <= 16'hFFFF;
rommem[7821] <= 16'hFFFF;
rommem[7822] <= 16'hFFFF;
rommem[7823] <= 16'hFFFF;
rommem[7824] <= 16'hFFFF;
rommem[7825] <= 16'hFFFF;
rommem[7826] <= 16'hFFFF;
rommem[7827] <= 16'hFFFF;
rommem[7828] <= 16'hFFFF;
rommem[7829] <= 16'hFFFF;
rommem[7830] <= 16'hFFFF;
rommem[7831] <= 16'hFFFF;
rommem[7832] <= 16'hFFFF;
rommem[7833] <= 16'hFFFF;
rommem[7834] <= 16'hFFFF;
rommem[7835] <= 16'hFFFF;
rommem[7836] <= 16'hFFFF;
rommem[7837] <= 16'hFFFF;
rommem[7838] <= 16'hFFFF;
rommem[7839] <= 16'hFFFF;
rommem[7840] <= 16'hFFFF;
rommem[7841] <= 16'hFFFF;
rommem[7842] <= 16'hFFFF;
rommem[7843] <= 16'hFFFF;
rommem[7844] <= 16'hFFFF;
rommem[7845] <= 16'hFFFF;
rommem[7846] <= 16'hFFFF;
rommem[7847] <= 16'hFFFF;
rommem[7848] <= 16'hFFFF;
rommem[7849] <= 16'hFFFF;
rommem[7850] <= 16'hFFFF;
rommem[7851] <= 16'hFFFF;
rommem[7852] <= 16'hFFFF;
rommem[7853] <= 16'hFFFF;
rommem[7854] <= 16'hFFFF;
rommem[7855] <= 16'hFFFF;
rommem[7856] <= 16'hFFFF;
rommem[7857] <= 16'hFFFF;
rommem[7858] <= 16'hFFFF;
rommem[7859] <= 16'hFFFF;
rommem[7860] <= 16'hFFFF;
rommem[7861] <= 16'hFFFF;
rommem[7862] <= 16'hFFFF;
rommem[7863] <= 16'hFFFF;
rommem[7864] <= 16'hFFFF;
rommem[7865] <= 16'hFFFF;
rommem[7866] <= 16'hFFFF;
rommem[7867] <= 16'hFFFF;
rommem[7868] <= 16'hFFFF;
rommem[7869] <= 16'hFFFF;
rommem[7870] <= 16'hFFFF;
rommem[7871] <= 16'hFFFF;
rommem[7872] <= 16'hFFFF;
rommem[7873] <= 16'hFFFF;
rommem[7874] <= 16'hFFFF;
rommem[7875] <= 16'hFFFF;
rommem[7876] <= 16'hFFFF;
rommem[7877] <= 16'hFFFF;
rommem[7878] <= 16'hFFFF;
rommem[7879] <= 16'hFFFF;
rommem[7880] <= 16'hFFFF;
rommem[7881] <= 16'hFFFF;
rommem[7882] <= 16'hFFFF;
rommem[7883] <= 16'hFFFF;
rommem[7884] <= 16'hFFFF;
rommem[7885] <= 16'hFFFF;
rommem[7886] <= 16'hFFFF;
rommem[7887] <= 16'hFFFF;
rommem[7888] <= 16'hFFFF;
rommem[7889] <= 16'hFFFF;
rommem[7890] <= 16'hFFFF;
rommem[7891] <= 16'hFFFF;
rommem[7892] <= 16'hFFFF;
rommem[7893] <= 16'hFFFF;
rommem[7894] <= 16'hFFFF;
rommem[7895] <= 16'hFFFF;
rommem[7896] <= 16'hFFFF;
rommem[7897] <= 16'hFFFF;
rommem[7898] <= 16'hFFFF;
rommem[7899] <= 16'hFFFF;
rommem[7900] <= 16'hFFFF;
rommem[7901] <= 16'hFFFF;
rommem[7902] <= 16'hFFFF;
rommem[7903] <= 16'hFFFF;
rommem[7904] <= 16'hFFFF;
rommem[7905] <= 16'hFFFF;
rommem[7906] <= 16'hFFFF;
rommem[7907] <= 16'hFFFF;
rommem[7908] <= 16'hFFFF;
rommem[7909] <= 16'hFFFF;
rommem[7910] <= 16'hFFFF;
rommem[7911] <= 16'hFFFF;
rommem[7912] <= 16'hFFFF;
rommem[7913] <= 16'hFFFF;
rommem[7914] <= 16'hFFFF;
rommem[7915] <= 16'hFFFF;
rommem[7916] <= 16'hFFFF;
rommem[7917] <= 16'hFFFF;
rommem[7918] <= 16'hFFFF;
rommem[7919] <= 16'hFFFF;
rommem[7920] <= 16'hFFFF;
rommem[7921] <= 16'hFFFF;
rommem[7922] <= 16'hFFFF;
rommem[7923] <= 16'hFFFF;
rommem[7924] <= 16'hFFFF;
rommem[7925] <= 16'hFFFF;
rommem[7926] <= 16'hFFFF;
rommem[7927] <= 16'hFFFF;
rommem[7928] <= 16'hFFFF;
rommem[7929] <= 16'hFFFF;
rommem[7930] <= 16'hFFFF;
rommem[7931] <= 16'hFFFF;
rommem[7932] <= 16'hFFFF;
rommem[7933] <= 16'hFFFF;
rommem[7934] <= 16'hFFFF;
rommem[7935] <= 16'hFFFF;
rommem[7936] <= 16'hFFFF;
rommem[7937] <= 16'hFFFF;
rommem[7938] <= 16'hFFFF;
rommem[7939] <= 16'hFFFF;
rommem[7940] <= 16'hFFFF;
rommem[7941] <= 16'hFFFF;
rommem[7942] <= 16'hFFFF;
rommem[7943] <= 16'hFFFF;
rommem[7944] <= 16'hFFFF;
rommem[7945] <= 16'hFFFF;
rommem[7946] <= 16'hFFFF;
rommem[7947] <= 16'hFFFF;
rommem[7948] <= 16'hFFFF;
rommem[7949] <= 16'hFFFF;
rommem[7950] <= 16'hFFFF;
rommem[7951] <= 16'hFFFF;
rommem[7952] <= 16'hFFFF;
rommem[7953] <= 16'hFFFF;
rommem[7954] <= 16'hFFFF;
rommem[7955] <= 16'hFFFF;
rommem[7956] <= 16'hFFFF;
rommem[7957] <= 16'hFFFF;
rommem[7958] <= 16'hFFFF;
rommem[7959] <= 16'hFFFF;
rommem[7960] <= 16'hFFFF;
rommem[7961] <= 16'hFFFF;
rommem[7962] <= 16'hFFFF;
rommem[7963] <= 16'hFFFF;
rommem[7964] <= 16'hFFFF;
rommem[7965] <= 16'hFFFF;
rommem[7966] <= 16'hFFFF;
rommem[7967] <= 16'hFFFF;
rommem[7968] <= 16'hFFFF;
rommem[7969] <= 16'hFFFF;
rommem[7970] <= 16'hFFFF;
rommem[7971] <= 16'hFFFF;
rommem[7972] <= 16'hFFFF;
rommem[7973] <= 16'hFFFF;
rommem[7974] <= 16'hFFFF;
rommem[7975] <= 16'hFFFF;
rommem[7976] <= 16'hFFFF;
rommem[7977] <= 16'hFFFF;
rommem[7978] <= 16'hFFFF;
rommem[7979] <= 16'hFFFF;
rommem[7980] <= 16'hFFFF;
rommem[7981] <= 16'hFFFF;
rommem[7982] <= 16'hFFFF;
rommem[7983] <= 16'hFFFF;
rommem[7984] <= 16'hFFFF;
rommem[7985] <= 16'hFFFF;
rommem[7986] <= 16'hFFFF;
rommem[7987] <= 16'hFFFF;
rommem[7988] <= 16'hFFFF;
rommem[7989] <= 16'hFFFF;
rommem[7990] <= 16'hFFFF;
rommem[7991] <= 16'hFFFF;
rommem[7992] <= 16'hFFFF;
rommem[7993] <= 16'hFFFF;
rommem[7994] <= 16'hFFFF;
rommem[7995] <= 16'hFFFF;
rommem[7996] <= 16'hFFFF;
rommem[7997] <= 16'hFFFF;
rommem[7998] <= 16'hFFFF;
rommem[7999] <= 16'hFFFF;
rommem[8000] <= 16'hFFFF;
rommem[8001] <= 16'hFFFF;
rommem[8002] <= 16'hFFFF;
rommem[8003] <= 16'hFFFF;
rommem[8004] <= 16'hFFFF;
rommem[8005] <= 16'hFFFF;
rommem[8006] <= 16'hFFFF;
rommem[8007] <= 16'hFFFF;
rommem[8008] <= 16'hFFFF;
rommem[8009] <= 16'hFFFF;
rommem[8010] <= 16'hFFFF;
rommem[8011] <= 16'hFFFF;
rommem[8012] <= 16'hFFFF;
rommem[8013] <= 16'hFFFF;
rommem[8014] <= 16'hFFFF;
rommem[8015] <= 16'hFFFF;
rommem[8016] <= 16'hFFFF;
rommem[8017] <= 16'hFFFF;
rommem[8018] <= 16'hFFFF;
rommem[8019] <= 16'hFFFF;
rommem[8020] <= 16'hFFFF;
rommem[8021] <= 16'hFFFF;
rommem[8022] <= 16'hFFFF;
rommem[8023] <= 16'hFFFF;
rommem[8024] <= 16'hFFFF;
rommem[8025] <= 16'hFFFF;
rommem[8026] <= 16'hFFFF;
rommem[8027] <= 16'hFFFF;
rommem[8028] <= 16'hFFFF;
rommem[8029] <= 16'hFFFF;
rommem[8030] <= 16'hFFFF;
rommem[8031] <= 16'hFFFF;
rommem[8032] <= 16'hFFFF;
rommem[8033] <= 16'hFFFF;
rommem[8034] <= 16'hFFFF;
rommem[8035] <= 16'hFFFF;
rommem[8036] <= 16'hFFFF;
rommem[8037] <= 16'hFFFF;
rommem[8038] <= 16'hFFFF;
rommem[8039] <= 16'hFFFF;
rommem[8040] <= 16'hFFFF;
rommem[8041] <= 16'hFFFF;
rommem[8042] <= 16'hFFFF;
rommem[8043] <= 16'hFFFF;
rommem[8044] <= 16'hFFFF;
rommem[8045] <= 16'hFFFF;
rommem[8046] <= 16'hFFFF;
rommem[8047] <= 16'hFFFF;
rommem[8048] <= 16'hFFFF;
rommem[8049] <= 16'hFFFF;
rommem[8050] <= 16'hFFFF;
rommem[8051] <= 16'hFFFF;
rommem[8052] <= 16'hFFFF;
rommem[8053] <= 16'hFFFF;
rommem[8054] <= 16'hFFFF;
rommem[8055] <= 16'hFFFF;
rommem[8056] <= 16'hFFFF;
rommem[8057] <= 16'hFFFF;
rommem[8058] <= 16'hFFFF;
rommem[8059] <= 16'hFFFF;
rommem[8060] <= 16'hFFFF;
rommem[8061] <= 16'hFFFF;
rommem[8062] <= 16'hFFFF;
rommem[8063] <= 16'hFFFF;
rommem[8064] <= 16'hFFFF;
rommem[8065] <= 16'hFFFF;
rommem[8066] <= 16'hFFFF;
rommem[8067] <= 16'hFFFF;
rommem[8068] <= 16'hFFFF;
rommem[8069] <= 16'hFFFF;
rommem[8070] <= 16'hFFFF;
rommem[8071] <= 16'hFFFF;
rommem[8072] <= 16'hFFFF;
rommem[8073] <= 16'hFFFF;
rommem[8074] <= 16'hFFFF;
rommem[8075] <= 16'hFFFF;
rommem[8076] <= 16'hFFFF;
rommem[8077] <= 16'hFFFF;
rommem[8078] <= 16'hFFFF;
rommem[8079] <= 16'hFFFF;
rommem[8080] <= 16'hFFFF;
rommem[8081] <= 16'hFFFF;
rommem[8082] <= 16'hFFFF;
rommem[8083] <= 16'hFFFF;
rommem[8084] <= 16'hFFFF;
rommem[8085] <= 16'hFFFF;
rommem[8086] <= 16'hFFFF;
rommem[8087] <= 16'hFFFF;
rommem[8088] <= 16'hFFFF;
rommem[8089] <= 16'hFFFF;
rommem[8090] <= 16'hFFFF;
rommem[8091] <= 16'hFFFF;
rommem[8092] <= 16'hFFFF;
rommem[8093] <= 16'hFFFF;
rommem[8094] <= 16'hFFFF;
rommem[8095] <= 16'hFFFF;
rommem[8096] <= 16'hFFFF;
rommem[8097] <= 16'hFFFF;
rommem[8098] <= 16'hFFFF;
rommem[8099] <= 16'hFFFF;
rommem[8100] <= 16'hFFFF;
rommem[8101] <= 16'hFFFF;
rommem[8102] <= 16'hFFFF;
rommem[8103] <= 16'hFFFF;
rommem[8104] <= 16'hFFFF;
rommem[8105] <= 16'hFFFF;
rommem[8106] <= 16'hFFFF;
rommem[8107] <= 16'hFFFF;
rommem[8108] <= 16'hFFFF;
rommem[8109] <= 16'hFFFF;
rommem[8110] <= 16'hFFFF;
rommem[8111] <= 16'hFFFF;
rommem[8112] <= 16'hFFFF;
rommem[8113] <= 16'hFFFF;
rommem[8114] <= 16'hFFFF;
rommem[8115] <= 16'hFFFF;
rommem[8116] <= 16'hFFFF;
rommem[8117] <= 16'hFFFF;
rommem[8118] <= 16'hFFFF;
rommem[8119] <= 16'hFFFF;
rommem[8120] <= 16'hFFFF;
rommem[8121] <= 16'hFFFF;
rommem[8122] <= 16'hFFFF;
rommem[8123] <= 16'hFFFF;
rommem[8124] <= 16'hFFFF;
rommem[8125] <= 16'hFFFF;
rommem[8126] <= 16'hFFFF;
rommem[8127] <= 16'hFFFF;
rommem[8128] <= 16'hFFFF;
rommem[8129] <= 16'hFFFF;
rommem[8130] <= 16'hFFFF;
rommem[8131] <= 16'hFFFF;
rommem[8132] <= 16'hFFFF;
rommem[8133] <= 16'hFFFF;
rommem[8134] <= 16'hFFFF;
rommem[8135] <= 16'hFFFF;
rommem[8136] <= 16'hFFFF;
rommem[8137] <= 16'hFFFF;
rommem[8138] <= 16'hFFFF;
rommem[8139] <= 16'hFFFF;
rommem[8140] <= 16'hFFFF;
rommem[8141] <= 16'hFFFF;
rommem[8142] <= 16'hFFFF;
rommem[8143] <= 16'hFFFF;
rommem[8144] <= 16'hFFFF;
rommem[8145] <= 16'hFFFF;
rommem[8146] <= 16'hFFFF;
rommem[8147] <= 16'hFFFF;
rommem[8148] <= 16'hFFFF;
rommem[8149] <= 16'hFFFF;
rommem[8150] <= 16'hFFFF;
rommem[8151] <= 16'hFFFF;
rommem[8152] <= 16'hFFFF;
rommem[8153] <= 16'hFFFF;
rommem[8154] <= 16'hFFFF;
rommem[8155] <= 16'hFFFF;
rommem[8156] <= 16'hFFFF;
rommem[8157] <= 16'hFFFF;
rommem[8158] <= 16'hFFFF;
rommem[8159] <= 16'hFFFF;
rommem[8160] <= 16'hFFFF;
rommem[8161] <= 16'hFFFF;
rommem[8162] <= 16'hFFFF;
rommem[8163] <= 16'hFFFF;
rommem[8164] <= 16'hFFFF;
rommem[8165] <= 16'hFFFF;
rommem[8166] <= 16'hFFFF;
rommem[8167] <= 16'hFFFF;
rommem[8168] <= 16'hFFFF;
rommem[8169] <= 16'hFFFF;
rommem[8170] <= 16'hFFFF;
rommem[8171] <= 16'hFFFF;
rommem[8172] <= 16'hFFFF;
rommem[8173] <= 16'hFFFF;
rommem[8174] <= 16'hFFFF;
rommem[8175] <= 16'hFFFF;
rommem[8176] <= 16'hFFFF;
rommem[8177] <= 16'hFFFF;
rommem[8178] <= 16'hFFFF;
rommem[8179] <= 16'hFFFF;
rommem[8180] <= 16'hFFFF;
rommem[8181] <= 16'hFFFF;
rommem[8182] <= 16'hFFFF;
rommem[8183] <= 16'hFFFF;
rommem[8184] <= 16'hFFFF;
rommem[8185] <= 16'hFFFF;
rommem[8186] <= 16'hFFFF;
rommem[8187] <= 16'hFFFF;
rommem[8188] <= 16'hFFFF;
rommem[8189] <= 16'hFFFF;
rommem[8190] <= 16'hFFFF;
rommem[8191] <= 16'hFFFF;
rommem[8192] <= 16'hFFFF;
rommem[8193] <= 16'hFFFF;
rommem[8194] <= 16'hFFFF;
rommem[8195] <= 16'hFFFF;
rommem[8196] <= 16'hFFFF;
rommem[8197] <= 16'hFFFF;
rommem[8198] <= 16'hFFFF;
rommem[8199] <= 16'hFFFF;
rommem[8200] <= 16'hFFFF;
rommem[8201] <= 16'hFFFF;
rommem[8202] <= 16'hFFFF;
rommem[8203] <= 16'hFFFF;
rommem[8204] <= 16'hFFFF;
rommem[8205] <= 16'hFFFF;
rommem[8206] <= 16'hFFFF;
rommem[8207] <= 16'hFFFF;
rommem[8208] <= 16'hFFFF;
rommem[8209] <= 16'hFFFF;
rommem[8210] <= 16'hFFFF;
rommem[8211] <= 16'hFFFF;
rommem[8212] <= 16'hFFFF;
rommem[8213] <= 16'hFFFF;
rommem[8214] <= 16'hFFFF;
rommem[8215] <= 16'hFFFF;
rommem[8216] <= 16'hFFFF;
rommem[8217] <= 16'hFFFF;
rommem[8218] <= 16'hFFFF;
rommem[8219] <= 16'hFFFF;
rommem[8220] <= 16'hFFFF;
rommem[8221] <= 16'hFFFF;
rommem[8222] <= 16'hFFFF;
rommem[8223] <= 16'hFFFF;
rommem[8224] <= 16'hFFFF;
rommem[8225] <= 16'hFFFF;
rommem[8226] <= 16'hFFFF;
rommem[8227] <= 16'hFFFF;
rommem[8228] <= 16'hFFFF;
rommem[8229] <= 16'hFFFF;
rommem[8230] <= 16'hFFFF;
rommem[8231] <= 16'hFFFF;
rommem[8232] <= 16'hFFFF;
rommem[8233] <= 16'hFFFF;
rommem[8234] <= 16'hFFFF;
rommem[8235] <= 16'hFFFF;
rommem[8236] <= 16'hFFFF;
rommem[8237] <= 16'hFFFF;
rommem[8238] <= 16'hFFFF;
rommem[8239] <= 16'hFFFF;
rommem[8240] <= 16'hFFFF;
rommem[8241] <= 16'hFFFF;
rommem[8242] <= 16'hFFFF;
rommem[8243] <= 16'hFFFF;
rommem[8244] <= 16'hFFFF;
rommem[8245] <= 16'hFFFF;
rommem[8246] <= 16'hFFFF;
rommem[8247] <= 16'hFFFF;
rommem[8248] <= 16'hFFFF;
rommem[8249] <= 16'hFFFF;
rommem[8250] <= 16'hFFFF;
rommem[8251] <= 16'hFFFF;
rommem[8252] <= 16'hFFFF;
rommem[8253] <= 16'hFFFF;
rommem[8254] <= 16'hFFFF;
rommem[8255] <= 16'hFFFF;
rommem[8256] <= 16'hFFFF;
rommem[8257] <= 16'hFFFF;
rommem[8258] <= 16'hFFFF;
rommem[8259] <= 16'hFFFF;
rommem[8260] <= 16'hFFFF;
rommem[8261] <= 16'hFFFF;
rommem[8262] <= 16'hFFFF;
rommem[8263] <= 16'hFFFF;
rommem[8264] <= 16'hFFFF;
rommem[8265] <= 16'hFFFF;
rommem[8266] <= 16'hFFFF;
rommem[8267] <= 16'hFFFF;
rommem[8268] <= 16'hFFFF;
rommem[8269] <= 16'hFFFF;
rommem[8270] <= 16'hFFFF;
rommem[8271] <= 16'hFFFF;
rommem[8272] <= 16'hFFFF;
rommem[8273] <= 16'hFFFF;
rommem[8274] <= 16'hFFFF;
rommem[8275] <= 16'hFFFF;
rommem[8276] <= 16'hFFFF;
rommem[8277] <= 16'hFFFF;
rommem[8278] <= 16'hFFFF;
rommem[8279] <= 16'hFFFF;
rommem[8280] <= 16'hFFFF;
rommem[8281] <= 16'hFFFF;
rommem[8282] <= 16'hFFFF;
rommem[8283] <= 16'hFFFF;
rommem[8284] <= 16'hFFFF;
rommem[8285] <= 16'hFFFF;
rommem[8286] <= 16'hFFFF;
rommem[8287] <= 16'hFFFF;
rommem[8288] <= 16'hFFFF;
rommem[8289] <= 16'hFFFF;
rommem[8290] <= 16'hFFFF;
rommem[8291] <= 16'hFFFF;
rommem[8292] <= 16'hFFFF;
rommem[8293] <= 16'hFFFF;
rommem[8294] <= 16'hFFFF;
rommem[8295] <= 16'hFFFF;
rommem[8296] <= 16'hFFFF;
rommem[8297] <= 16'hFFFF;
rommem[8298] <= 16'hFFFF;
rommem[8299] <= 16'hFFFF;
rommem[8300] <= 16'hFFFF;
rommem[8301] <= 16'hFFFF;
rommem[8302] <= 16'hFFFF;
rommem[8303] <= 16'hFFFF;
rommem[8304] <= 16'hFFFF;
rommem[8305] <= 16'hFFFF;
rommem[8306] <= 16'hFFFF;
rommem[8307] <= 16'hFFFF;
rommem[8308] <= 16'hFFFF;
rommem[8309] <= 16'hFFFF;
rommem[8310] <= 16'hFFFF;
rommem[8311] <= 16'hFFFF;
rommem[8312] <= 16'hFFFF;
rommem[8313] <= 16'hFFFF;
rommem[8314] <= 16'hFFFF;
rommem[8315] <= 16'hFFFF;
rommem[8316] <= 16'hFFFF;
rommem[8317] <= 16'hFFFF;
rommem[8318] <= 16'hFFFF;
rommem[8319] <= 16'hFFFF;
rommem[8320] <= 16'hFFFF;
rommem[8321] <= 16'hFFFF;
rommem[8322] <= 16'hFFFF;
rommem[8323] <= 16'hFFFF;
rommem[8324] <= 16'hFFFF;
rommem[8325] <= 16'hFFFF;
rommem[8326] <= 16'hFFFF;
rommem[8327] <= 16'hFFFF;
rommem[8328] <= 16'hFFFF;
rommem[8329] <= 16'hFFFF;
rommem[8330] <= 16'hFFFF;
rommem[8331] <= 16'hFFFF;
rommem[8332] <= 16'hFFFF;
rommem[8333] <= 16'hFFFF;
rommem[8334] <= 16'hFFFF;
rommem[8335] <= 16'hFFFF;
rommem[8336] <= 16'hFFFF;
rommem[8337] <= 16'hFFFF;
rommem[8338] <= 16'hFFFF;
rommem[8339] <= 16'hFFFF;
rommem[8340] <= 16'hFFFF;
rommem[8341] <= 16'hFFFF;
rommem[8342] <= 16'hFFFF;
rommem[8343] <= 16'hFFFF;
rommem[8344] <= 16'hFFFF;
rommem[8345] <= 16'hFFFF;
rommem[8346] <= 16'hFFFF;
rommem[8347] <= 16'hFFFF;
rommem[8348] <= 16'hFFFF;
rommem[8349] <= 16'hFFFF;
rommem[8350] <= 16'hFFFF;
rommem[8351] <= 16'hFFFF;
rommem[8352] <= 16'hFFFF;
rommem[8353] <= 16'hFFFF;
rommem[8354] <= 16'hFFFF;
rommem[8355] <= 16'hFFFF;
rommem[8356] <= 16'hFFFF;
rommem[8357] <= 16'hFFFF;
rommem[8358] <= 16'hFFFF;
rommem[8359] <= 16'hFFFF;
rommem[8360] <= 16'hFFFF;
rommem[8361] <= 16'hFFFF;
rommem[8362] <= 16'hFFFF;
rommem[8363] <= 16'hFFFF;
rommem[8364] <= 16'hFFFF;
rommem[8365] <= 16'hFFFF;
rommem[8366] <= 16'hFFFF;
rommem[8367] <= 16'hFFFF;
rommem[8368] <= 16'hFFFF;
rommem[8369] <= 16'hFFFF;
rommem[8370] <= 16'hFFFF;
rommem[8371] <= 16'hFFFF;
rommem[8372] <= 16'hFFFF;
rommem[8373] <= 16'hFFFF;
rommem[8374] <= 16'hFFFF;
rommem[8375] <= 16'hFFFF;
rommem[8376] <= 16'hFFFF;
rommem[8377] <= 16'hFFFF;
rommem[8378] <= 16'hFFFF;
rommem[8379] <= 16'hFFFF;
rommem[8380] <= 16'hFFFF;
rommem[8381] <= 16'hFFFF;
rommem[8382] <= 16'hFFFF;
rommem[8383] <= 16'hFFFF;
rommem[8384] <= 16'hFFFF;
rommem[8385] <= 16'hFFFF;
rommem[8386] <= 16'hFFFF;
rommem[8387] <= 16'hFFFF;
rommem[8388] <= 16'hFFFF;
rommem[8389] <= 16'hFFFF;
rommem[8390] <= 16'hFFFF;
rommem[8391] <= 16'hFFFF;
rommem[8392] <= 16'hFFFF;
rommem[8393] <= 16'hFFFF;
rommem[8394] <= 16'hFFFF;
rommem[8395] <= 16'hFFFF;
rommem[8396] <= 16'hFFFF;
rommem[8397] <= 16'hFFFF;
rommem[8398] <= 16'hFFFF;
rommem[8399] <= 16'hFFFF;
rommem[8400] <= 16'hFFFF;
rommem[8401] <= 16'hFFFF;
rommem[8402] <= 16'hFFFF;
rommem[8403] <= 16'hFFFF;
rommem[8404] <= 16'hFFFF;
rommem[8405] <= 16'hFFFF;
rommem[8406] <= 16'hFFFF;
rommem[8407] <= 16'hFFFF;
rommem[8408] <= 16'hFFFF;
rommem[8409] <= 16'hFFFF;
rommem[8410] <= 16'hFFFF;
rommem[8411] <= 16'hFFFF;
rommem[8412] <= 16'hFFFF;
rommem[8413] <= 16'hFFFF;
rommem[8414] <= 16'hFFFF;
rommem[8415] <= 16'hFFFF;
rommem[8416] <= 16'hFFFF;
rommem[8417] <= 16'hFFFF;
rommem[8418] <= 16'hFFFF;
rommem[8419] <= 16'hFFFF;
rommem[8420] <= 16'hFFFF;
rommem[8421] <= 16'hFFFF;
rommem[8422] <= 16'hFFFF;
rommem[8423] <= 16'hFFFF;
rommem[8424] <= 16'hFFFF;
rommem[8425] <= 16'hFFFF;
rommem[8426] <= 16'hFFFF;
rommem[8427] <= 16'hFFFF;
rommem[8428] <= 16'hFFFF;
rommem[8429] <= 16'hFFFF;
rommem[8430] <= 16'hFFFF;
rommem[8431] <= 16'hFFFF;
rommem[8432] <= 16'hFFFF;
rommem[8433] <= 16'hFFFF;
rommem[8434] <= 16'hFFFF;
rommem[8435] <= 16'hFFFF;
rommem[8436] <= 16'hFFFF;
rommem[8437] <= 16'hFFFF;
rommem[8438] <= 16'hFFFF;
rommem[8439] <= 16'hFFFF;
rommem[8440] <= 16'hFFFF;
rommem[8441] <= 16'hFFFF;
rommem[8442] <= 16'hFFFF;
rommem[8443] <= 16'hFFFF;
rommem[8444] <= 16'hFFFF;
rommem[8445] <= 16'hFFFF;
rommem[8446] <= 16'hFFFF;
rommem[8447] <= 16'hFFFF;
rommem[8448] <= 16'hFFFF;
rommem[8449] <= 16'hFFFF;
rommem[8450] <= 16'hFFFF;
rommem[8451] <= 16'hFFFF;
rommem[8452] <= 16'hFFFF;
rommem[8453] <= 16'hFFFF;
rommem[8454] <= 16'hFFFF;
rommem[8455] <= 16'hFFFF;
rommem[8456] <= 16'hFFFF;
rommem[8457] <= 16'hFFFF;
rommem[8458] <= 16'hFFFF;
rommem[8459] <= 16'hFFFF;
rommem[8460] <= 16'hFFFF;
rommem[8461] <= 16'hFFFF;
rommem[8462] <= 16'hFFFF;
rommem[8463] <= 16'hFFFF;
rommem[8464] <= 16'hFFFF;
rommem[8465] <= 16'hFFFF;
rommem[8466] <= 16'hFFFF;
rommem[8467] <= 16'hFFFF;
rommem[8468] <= 16'hFFFF;
rommem[8469] <= 16'hFFFF;
rommem[8470] <= 16'hFFFF;
rommem[8471] <= 16'hFFFF;
rommem[8472] <= 16'hFFFF;
rommem[8473] <= 16'hFFFF;
rommem[8474] <= 16'hFFFF;
rommem[8475] <= 16'hFFFF;
rommem[8476] <= 16'hFFFF;
rommem[8477] <= 16'hFFFF;
rommem[8478] <= 16'hFFFF;
rommem[8479] <= 16'hFFFF;
rommem[8480] <= 16'hFFFF;
rommem[8481] <= 16'hFFFF;
rommem[8482] <= 16'hFFFF;
rommem[8483] <= 16'hFFFF;
rommem[8484] <= 16'hFFFF;
rommem[8485] <= 16'hFFFF;
rommem[8486] <= 16'hFFFF;
rommem[8487] <= 16'hFFFF;
rommem[8488] <= 16'hFFFF;
rommem[8489] <= 16'hFFFF;
rommem[8490] <= 16'hFFFF;
rommem[8491] <= 16'hFFFF;
rommem[8492] <= 16'hFFFF;
rommem[8493] <= 16'hFFFF;
rommem[8494] <= 16'hFFFF;
rommem[8495] <= 16'hFFFF;
rommem[8496] <= 16'hFFFF;
rommem[8497] <= 16'hFFFF;
rommem[8498] <= 16'hFFFF;
rommem[8499] <= 16'hFFFF;
rommem[8500] <= 16'hFFFF;
rommem[8501] <= 16'hFFFF;
rommem[8502] <= 16'hFFFF;
rommem[8503] <= 16'hFFFF;
rommem[8504] <= 16'hFFFF;
rommem[8505] <= 16'hFFFF;
rommem[8506] <= 16'hFFFF;
rommem[8507] <= 16'hFFFF;
rommem[8508] <= 16'hFFFF;
rommem[8509] <= 16'hFFFF;
rommem[8510] <= 16'hFFFF;
rommem[8511] <= 16'hFFFF;
rommem[8512] <= 16'hFFFF;
rommem[8513] <= 16'hFFFF;
rommem[8514] <= 16'hFFFF;
rommem[8515] <= 16'hFFFF;
rommem[8516] <= 16'hFFFF;
rommem[8517] <= 16'hFFFF;
rommem[8518] <= 16'hFFFF;
rommem[8519] <= 16'hFFFF;
rommem[8520] <= 16'hFFFF;
rommem[8521] <= 16'hFFFF;
rommem[8522] <= 16'hFFFF;
rommem[8523] <= 16'hFFFF;
rommem[8524] <= 16'hFFFF;
rommem[8525] <= 16'hFFFF;
rommem[8526] <= 16'hFFFF;
rommem[8527] <= 16'hFFFF;
rommem[8528] <= 16'hFFFF;
rommem[8529] <= 16'hFFFF;
rommem[8530] <= 16'hFFFF;
rommem[8531] <= 16'hFFFF;
rommem[8532] <= 16'hFFFF;
rommem[8533] <= 16'hFFFF;
rommem[8534] <= 16'hFFFF;
rommem[8535] <= 16'hFFFF;
rommem[8536] <= 16'hFFFF;
rommem[8537] <= 16'hFFFF;
rommem[8538] <= 16'hFFFF;
rommem[8539] <= 16'hFFFF;
rommem[8540] <= 16'hFFFF;
rommem[8541] <= 16'hFFFF;
rommem[8542] <= 16'hFFFF;
rommem[8543] <= 16'hFFFF;
rommem[8544] <= 16'hFFFF;
rommem[8545] <= 16'hFFFF;
rommem[8546] <= 16'hFFFF;
rommem[8547] <= 16'hFFFF;
rommem[8548] <= 16'hFFFF;
rommem[8549] <= 16'hFFFF;
rommem[8550] <= 16'hFFFF;
rommem[8551] <= 16'hFFFF;
rommem[8552] <= 16'hFFFF;
rommem[8553] <= 16'hFFFF;
rommem[8554] <= 16'hFFFF;
rommem[8555] <= 16'hFFFF;
rommem[8556] <= 16'hFFFF;
rommem[8557] <= 16'hFFFF;
rommem[8558] <= 16'hFFFF;
rommem[8559] <= 16'hFFFF;
rommem[8560] <= 16'hFFFF;
rommem[8561] <= 16'hFFFF;
rommem[8562] <= 16'hFFFF;
rommem[8563] <= 16'hFFFF;
rommem[8564] <= 16'hFFFF;
rommem[8565] <= 16'hFFFF;
rommem[8566] <= 16'hFFFF;
rommem[8567] <= 16'hFFFF;
rommem[8568] <= 16'hFFFF;
rommem[8569] <= 16'hFFFF;
rommem[8570] <= 16'hFFFF;
rommem[8571] <= 16'hFFFF;
rommem[8572] <= 16'hFFFF;
rommem[8573] <= 16'hFFFF;
rommem[8574] <= 16'hFFFF;
rommem[8575] <= 16'hFFFF;
rommem[8576] <= 16'hFFFF;
rommem[8577] <= 16'hFFFF;
rommem[8578] <= 16'hFFFF;
rommem[8579] <= 16'hFFFF;
rommem[8580] <= 16'hFFFF;
rommem[8581] <= 16'hFFFF;
rommem[8582] <= 16'hFFFF;
rommem[8583] <= 16'hFFFF;
rommem[8584] <= 16'hFFFF;
rommem[8585] <= 16'hFFFF;
rommem[8586] <= 16'hFFFF;
rommem[8587] <= 16'hFFFF;
rommem[8588] <= 16'hFFFF;
rommem[8589] <= 16'hFFFF;
rommem[8590] <= 16'hFFFF;
rommem[8591] <= 16'hFFFF;
rommem[8592] <= 16'hFFFF;
rommem[8593] <= 16'hFFFF;
rommem[8594] <= 16'hFFFF;
rommem[8595] <= 16'hFFFF;
rommem[8596] <= 16'hFFFF;
rommem[8597] <= 16'hFFFF;
rommem[8598] <= 16'hFFFF;
rommem[8599] <= 16'hFFFF;
rommem[8600] <= 16'hFFFF;
rommem[8601] <= 16'hFFFF;
rommem[8602] <= 16'hFFFF;
rommem[8603] <= 16'hFFFF;
rommem[8604] <= 16'hFFFF;
rommem[8605] <= 16'hFFFF;
rommem[8606] <= 16'hFFFF;
rommem[8607] <= 16'hFFFF;
rommem[8608] <= 16'hFFFF;
rommem[8609] <= 16'hFFFF;
rommem[8610] <= 16'hFFFF;
rommem[8611] <= 16'hFFFF;
rommem[8612] <= 16'hFFFF;
rommem[8613] <= 16'hFFFF;
rommem[8614] <= 16'hFFFF;
rommem[8615] <= 16'hFFFF;
rommem[8616] <= 16'hFFFF;
rommem[8617] <= 16'hFFFF;
rommem[8618] <= 16'hFFFF;
rommem[8619] <= 16'hFFFF;
rommem[8620] <= 16'hFFFF;
rommem[8621] <= 16'hFFFF;
rommem[8622] <= 16'hFFFF;
rommem[8623] <= 16'hFFFF;
rommem[8624] <= 16'hFFFF;
rommem[8625] <= 16'hFFFF;
rommem[8626] <= 16'hFFFF;
rommem[8627] <= 16'hFFFF;
rommem[8628] <= 16'hFFFF;
rommem[8629] <= 16'hFFFF;
rommem[8630] <= 16'hFFFF;
rommem[8631] <= 16'hFFFF;
rommem[8632] <= 16'hFFFF;
rommem[8633] <= 16'hFFFF;
rommem[8634] <= 16'hFFFF;
rommem[8635] <= 16'hFFFF;
rommem[8636] <= 16'hFFFF;
rommem[8637] <= 16'hFFFF;
rommem[8638] <= 16'hFFFF;
rommem[8639] <= 16'hFFFF;
rommem[8640] <= 16'hFFFF;
rommem[8641] <= 16'hFFFF;
rommem[8642] <= 16'hFFFF;
rommem[8643] <= 16'hFFFF;
rommem[8644] <= 16'hFFFF;
rommem[8645] <= 16'hFFFF;
rommem[8646] <= 16'hFFFF;
rommem[8647] <= 16'hFFFF;
rommem[8648] <= 16'hFFFF;
rommem[8649] <= 16'hFFFF;
rommem[8650] <= 16'hFFFF;
rommem[8651] <= 16'hFFFF;
rommem[8652] <= 16'hFFFF;
rommem[8653] <= 16'hFFFF;
rommem[8654] <= 16'hFFFF;
rommem[8655] <= 16'hFFFF;
rommem[8656] <= 16'hFFFF;
rommem[8657] <= 16'hFFFF;
rommem[8658] <= 16'hFFFF;
rommem[8659] <= 16'hFFFF;
rommem[8660] <= 16'hFFFF;
rommem[8661] <= 16'hFFFF;
rommem[8662] <= 16'hFFFF;
rommem[8663] <= 16'hFFFF;
rommem[8664] <= 16'hFFFF;
rommem[8665] <= 16'hFFFF;
rommem[8666] <= 16'hFFFF;
rommem[8667] <= 16'hFFFF;
rommem[8668] <= 16'hFFFF;
rommem[8669] <= 16'hFFFF;
rommem[8670] <= 16'hFFFF;
rommem[8671] <= 16'hFFFF;
rommem[8672] <= 16'hFFFF;
rommem[8673] <= 16'hFFFF;
rommem[8674] <= 16'hFFFF;
rommem[8675] <= 16'hFFFF;
rommem[8676] <= 16'hFFFF;
rommem[8677] <= 16'hFFFF;
rommem[8678] <= 16'hFFFF;
rommem[8679] <= 16'hFFFF;
rommem[8680] <= 16'hFFFF;
rommem[8681] <= 16'hFFFF;
rommem[8682] <= 16'hFFFF;
rommem[8683] <= 16'hFFFF;
rommem[8684] <= 16'hFFFF;
rommem[8685] <= 16'hFFFF;
rommem[8686] <= 16'hFFFF;
rommem[8687] <= 16'hFFFF;
rommem[8688] <= 16'hFFFF;
rommem[8689] <= 16'hFFFF;
rommem[8690] <= 16'hFFFF;
rommem[8691] <= 16'hFFFF;
rommem[8692] <= 16'hFFFF;
rommem[8693] <= 16'hFFFF;
rommem[8694] <= 16'hFFFF;
rommem[8695] <= 16'hFFFF;
rommem[8696] <= 16'hFFFF;
rommem[8697] <= 16'hFFFF;
rommem[8698] <= 16'hFFFF;
rommem[8699] <= 16'hFFFF;
rommem[8700] <= 16'hFFFF;
rommem[8701] <= 16'hFFFF;
rommem[8702] <= 16'hFFFF;
rommem[8703] <= 16'hFFFF;
rommem[8704] <= 16'hFFFF;
rommem[8705] <= 16'hFFFF;
rommem[8706] <= 16'hFFFF;
rommem[8707] <= 16'hFFFF;
rommem[8708] <= 16'hFFFF;
rommem[8709] <= 16'hFFFF;
rommem[8710] <= 16'hFFFF;
rommem[8711] <= 16'hFFFF;
rommem[8712] <= 16'hFFFF;
rommem[8713] <= 16'hFFFF;
rommem[8714] <= 16'hFFFF;
rommem[8715] <= 16'hFFFF;
rommem[8716] <= 16'hFFFF;
rommem[8717] <= 16'hFFFF;
rommem[8718] <= 16'hFFFF;
rommem[8719] <= 16'hFFFF;
rommem[8720] <= 16'hFFFF;
rommem[8721] <= 16'hFFFF;
rommem[8722] <= 16'hFFFF;
rommem[8723] <= 16'hFFFF;
rommem[8724] <= 16'hFFFF;
rommem[8725] <= 16'hFFFF;
rommem[8726] <= 16'hFFFF;
rommem[8727] <= 16'hFFFF;
rommem[8728] <= 16'hFFFF;
rommem[8729] <= 16'hFFFF;
rommem[8730] <= 16'hFFFF;
rommem[8731] <= 16'hFFFF;
rommem[8732] <= 16'hFFFF;
rommem[8733] <= 16'hFFFF;
rommem[8734] <= 16'hFFFF;
rommem[8735] <= 16'hFFFF;
rommem[8736] <= 16'hFFFF;
rommem[8737] <= 16'hFFFF;
rommem[8738] <= 16'hFFFF;
rommem[8739] <= 16'hFFFF;
rommem[8740] <= 16'hFFFF;
rommem[8741] <= 16'hFFFF;
rommem[8742] <= 16'hFFFF;
rommem[8743] <= 16'hFFFF;
rommem[8744] <= 16'hFFFF;
rommem[8745] <= 16'hFFFF;
rommem[8746] <= 16'hFFFF;
rommem[8747] <= 16'hFFFF;
rommem[8748] <= 16'hFFFF;
rommem[8749] <= 16'hFFFF;
rommem[8750] <= 16'hFFFF;
rommem[8751] <= 16'hFFFF;
rommem[8752] <= 16'hFFFF;
rommem[8753] <= 16'hFFFF;
rommem[8754] <= 16'hFFFF;
rommem[8755] <= 16'hFFFF;
rommem[8756] <= 16'hFFFF;
rommem[8757] <= 16'hFFFF;
rommem[8758] <= 16'hFFFF;
rommem[8759] <= 16'hFFFF;
rommem[8760] <= 16'hFFFF;
rommem[8761] <= 16'hFFFF;
rommem[8762] <= 16'hFFFF;
rommem[8763] <= 16'hFFFF;
rommem[8764] <= 16'hFFFF;
rommem[8765] <= 16'hFFFF;
rommem[8766] <= 16'hFFFF;
rommem[8767] <= 16'hFFFF;
rommem[8768] <= 16'hFFFF;
rommem[8769] <= 16'hFFFF;
rommem[8770] <= 16'hFFFF;
rommem[8771] <= 16'hFFFF;
rommem[8772] <= 16'hFFFF;
rommem[8773] <= 16'hFFFF;
rommem[8774] <= 16'hFFFF;
rommem[8775] <= 16'hFFFF;
rommem[8776] <= 16'hFFFF;
rommem[8777] <= 16'hFFFF;
rommem[8778] <= 16'hFFFF;
rommem[8779] <= 16'hFFFF;
rommem[8780] <= 16'hFFFF;
rommem[8781] <= 16'hFFFF;
rommem[8782] <= 16'hFFFF;
rommem[8783] <= 16'hFFFF;
rommem[8784] <= 16'hFFFF;
rommem[8785] <= 16'hFFFF;
rommem[8786] <= 16'hFFFF;
rommem[8787] <= 16'hFFFF;
rommem[8788] <= 16'hFFFF;
rommem[8789] <= 16'hFFFF;
rommem[8790] <= 16'hFFFF;
rommem[8791] <= 16'hFFFF;
rommem[8792] <= 16'hFFFF;
rommem[8793] <= 16'hFFFF;
rommem[8794] <= 16'hFFFF;
rommem[8795] <= 16'hFFFF;
rommem[8796] <= 16'hFFFF;
rommem[8797] <= 16'hFFFF;
rommem[8798] <= 16'hFFFF;
rommem[8799] <= 16'hFFFF;
rommem[8800] <= 16'hFFFF;
rommem[8801] <= 16'hFFFF;
rommem[8802] <= 16'hFFFF;
rommem[8803] <= 16'hFFFF;
rommem[8804] <= 16'hFFFF;
rommem[8805] <= 16'hFFFF;
rommem[8806] <= 16'hFFFF;
rommem[8807] <= 16'hFFFF;
rommem[8808] <= 16'hFFFF;
rommem[8809] <= 16'hFFFF;
rommem[8810] <= 16'hFFFF;
rommem[8811] <= 16'hFFFF;
rommem[8812] <= 16'hFFFF;
rommem[8813] <= 16'hFFFF;
rommem[8814] <= 16'hFFFF;
rommem[8815] <= 16'hFFFF;
rommem[8816] <= 16'hFFFF;
rommem[8817] <= 16'hFFFF;
rommem[8818] <= 16'hFFFF;
rommem[8819] <= 16'hFFFF;
rommem[8820] <= 16'hFFFF;
rommem[8821] <= 16'hFFFF;
rommem[8822] <= 16'hFFFF;
rommem[8823] <= 16'hFFFF;
rommem[8824] <= 16'hFFFF;
rommem[8825] <= 16'hFFFF;
rommem[8826] <= 16'hFFFF;
rommem[8827] <= 16'hFFFF;
rommem[8828] <= 16'hFFFF;
rommem[8829] <= 16'hFFFF;
rommem[8830] <= 16'hFFFF;
rommem[8831] <= 16'hFFFF;
rommem[8832] <= 16'hFFFF;
rommem[8833] <= 16'hFFFF;
rommem[8834] <= 16'hFFFF;
rommem[8835] <= 16'hFFFF;
rommem[8836] <= 16'hFFFF;
rommem[8837] <= 16'hFFFF;
rommem[8838] <= 16'hFFFF;
rommem[8839] <= 16'hFFFF;
rommem[8840] <= 16'hFFFF;
rommem[8841] <= 16'hFFFF;
rommem[8842] <= 16'hFFFF;
rommem[8843] <= 16'hFFFF;
rommem[8844] <= 16'hFFFF;
rommem[8845] <= 16'hFFFF;
rommem[8846] <= 16'hFFFF;
rommem[8847] <= 16'hFFFF;
rommem[8848] <= 16'hFFFF;
rommem[8849] <= 16'hFFFF;
rommem[8850] <= 16'hFFFF;
rommem[8851] <= 16'hFFFF;
rommem[8852] <= 16'hFFFF;
rommem[8853] <= 16'hFFFF;
rommem[8854] <= 16'hFFFF;
rommem[8855] <= 16'hFFFF;
rommem[8856] <= 16'hFFFF;
rommem[8857] <= 16'hFFFF;
rommem[8858] <= 16'hFFFF;
rommem[8859] <= 16'hFFFF;
rommem[8860] <= 16'hFFFF;
rommem[8861] <= 16'hFFFF;
rommem[8862] <= 16'hFFFF;
rommem[8863] <= 16'hFFFF;
rommem[8864] <= 16'hFFFF;
rommem[8865] <= 16'hFFFF;
rommem[8866] <= 16'hFFFF;
rommem[8867] <= 16'hFFFF;
rommem[8868] <= 16'hFFFF;
rommem[8869] <= 16'hFFFF;
rommem[8870] <= 16'hFFFF;
rommem[8871] <= 16'hFFFF;
rommem[8872] <= 16'hFFFF;
rommem[8873] <= 16'hFFFF;
rommem[8874] <= 16'hFFFF;
rommem[8875] <= 16'hFFFF;
rommem[8876] <= 16'hFFFF;
rommem[8877] <= 16'hFFFF;
rommem[8878] <= 16'hFFFF;
rommem[8879] <= 16'hFFFF;
rommem[8880] <= 16'hFFFF;
rommem[8881] <= 16'hFFFF;
rommem[8882] <= 16'hFFFF;
rommem[8883] <= 16'hFFFF;
rommem[8884] <= 16'hFFFF;
rommem[8885] <= 16'hFFFF;
rommem[8886] <= 16'hFFFF;
rommem[8887] <= 16'hFFFF;
rommem[8888] <= 16'hFFFF;
rommem[8889] <= 16'hFFFF;
rommem[8890] <= 16'hFFFF;
rommem[8891] <= 16'hFFFF;
rommem[8892] <= 16'hFFFF;
rommem[8893] <= 16'hFFFF;
rommem[8894] <= 16'hFFFF;
rommem[8895] <= 16'hFFFF;
rommem[8896] <= 16'hFFFF;
rommem[8897] <= 16'hFFFF;
rommem[8898] <= 16'hFFFF;
rommem[8899] <= 16'hFFFF;
rommem[8900] <= 16'hFFFF;
rommem[8901] <= 16'hFFFF;
rommem[8902] <= 16'hFFFF;
rommem[8903] <= 16'hFFFF;
rommem[8904] <= 16'hFFFF;
rommem[8905] <= 16'hFFFF;
rommem[8906] <= 16'hFFFF;
rommem[8907] <= 16'hFFFF;
rommem[8908] <= 16'hFFFF;
rommem[8909] <= 16'hFFFF;
rommem[8910] <= 16'hFFFF;
rommem[8911] <= 16'hFFFF;
rommem[8912] <= 16'hFFFF;
rommem[8913] <= 16'hFFFF;
rommem[8914] <= 16'hFFFF;
rommem[8915] <= 16'hFFFF;
rommem[8916] <= 16'hFFFF;
rommem[8917] <= 16'hFFFF;
rommem[8918] <= 16'hFFFF;
rommem[8919] <= 16'hFFFF;
rommem[8920] <= 16'hFFFF;
rommem[8921] <= 16'hFFFF;
rommem[8922] <= 16'hFFFF;
rommem[8923] <= 16'hFFFF;
rommem[8924] <= 16'hFFFF;
rommem[8925] <= 16'hFFFF;
rommem[8926] <= 16'hFFFF;
rommem[8927] <= 16'hFFFF;
rommem[8928] <= 16'hFFFF;
rommem[8929] <= 16'hFFFF;
rommem[8930] <= 16'hFFFF;
rommem[8931] <= 16'hFFFF;
rommem[8932] <= 16'hFFFF;
rommem[8933] <= 16'hFFFF;
rommem[8934] <= 16'hFFFF;
rommem[8935] <= 16'hFFFF;
rommem[8936] <= 16'hFFFF;
rommem[8937] <= 16'hFFFF;
rommem[8938] <= 16'hFFFF;
rommem[8939] <= 16'hFFFF;
rommem[8940] <= 16'hFFFF;
rommem[8941] <= 16'hFFFF;
rommem[8942] <= 16'hFFFF;
rommem[8943] <= 16'hFFFF;
rommem[8944] <= 16'hFFFF;
rommem[8945] <= 16'hFFFF;
rommem[8946] <= 16'hFFFF;
rommem[8947] <= 16'hFFFF;
rommem[8948] <= 16'hFFFF;
rommem[8949] <= 16'hFFFF;
rommem[8950] <= 16'hFFFF;
rommem[8951] <= 16'hFFFF;
rommem[8952] <= 16'hFFFF;
rommem[8953] <= 16'hFFFF;
rommem[8954] <= 16'hFFFF;
rommem[8955] <= 16'hFFFF;
rommem[8956] <= 16'hFFFF;
rommem[8957] <= 16'hFFFF;
rommem[8958] <= 16'hFFFF;
rommem[8959] <= 16'hFFFF;
rommem[8960] <= 16'hFFFF;
rommem[8961] <= 16'hFFFF;
rommem[8962] <= 16'hFFFF;
rommem[8963] <= 16'hFFFF;
rommem[8964] <= 16'hFFFF;
rommem[8965] <= 16'hFFFF;
rommem[8966] <= 16'hFFFF;
rommem[8967] <= 16'hFFFF;
rommem[8968] <= 16'hFFFF;
rommem[8969] <= 16'hFFFF;
rommem[8970] <= 16'hFFFF;
rommem[8971] <= 16'hFFFF;
rommem[8972] <= 16'hFFFF;
rommem[8973] <= 16'hFFFF;
rommem[8974] <= 16'hFFFF;
rommem[8975] <= 16'hFFFF;
rommem[8976] <= 16'hFFFF;
rommem[8977] <= 16'hFFFF;
rommem[8978] <= 16'hFFFF;
rommem[8979] <= 16'hFFFF;
rommem[8980] <= 16'hFFFF;
rommem[8981] <= 16'hFFFF;
rommem[8982] <= 16'hFFFF;
rommem[8983] <= 16'hFFFF;
rommem[8984] <= 16'hFFFF;
rommem[8985] <= 16'hFFFF;
rommem[8986] <= 16'hFFFF;
rommem[8987] <= 16'hFFFF;
rommem[8988] <= 16'hFFFF;
rommem[8989] <= 16'hFFFF;
rommem[8990] <= 16'hFFFF;
rommem[8991] <= 16'hFFFF;
rommem[8992] <= 16'hFFFF;
rommem[8993] <= 16'hFFFF;
rommem[8994] <= 16'hFFFF;
rommem[8995] <= 16'hFFFF;
rommem[8996] <= 16'hFFFF;
rommem[8997] <= 16'hFFFF;
rommem[8998] <= 16'hFFFF;
rommem[8999] <= 16'hFFFF;
rommem[9000] <= 16'hFFFF;
rommem[9001] <= 16'hFFFF;
rommem[9002] <= 16'hFFFF;
rommem[9003] <= 16'hFFFF;
rommem[9004] <= 16'hFFFF;
rommem[9005] <= 16'hFFFF;
rommem[9006] <= 16'hFFFF;
rommem[9007] <= 16'hFFFF;
rommem[9008] <= 16'hFFFF;
rommem[9009] <= 16'hFFFF;
rommem[9010] <= 16'hFFFF;
rommem[9011] <= 16'hFFFF;
rommem[9012] <= 16'hFFFF;
rommem[9013] <= 16'hFFFF;
rommem[9014] <= 16'hFFFF;
rommem[9015] <= 16'hFFFF;
rommem[9016] <= 16'hFFFF;
rommem[9017] <= 16'hFFFF;
rommem[9018] <= 16'hFFFF;
rommem[9019] <= 16'hFFFF;
rommem[9020] <= 16'hFFFF;
rommem[9021] <= 16'hFFFF;
rommem[9022] <= 16'hFFFF;
rommem[9023] <= 16'hFFFF;
rommem[9024] <= 16'hFFFF;
rommem[9025] <= 16'hFFFF;
rommem[9026] <= 16'hFFFF;
rommem[9027] <= 16'hFFFF;
rommem[9028] <= 16'hFFFF;
rommem[9029] <= 16'hFFFF;
rommem[9030] <= 16'hFFFF;
rommem[9031] <= 16'hFFFF;
rommem[9032] <= 16'hFFFF;
rommem[9033] <= 16'hFFFF;
rommem[9034] <= 16'hFFFF;
rommem[9035] <= 16'hFFFF;
rommem[9036] <= 16'hFFFF;
rommem[9037] <= 16'hFFFF;
rommem[9038] <= 16'hFFFF;
rommem[9039] <= 16'hFFFF;
rommem[9040] <= 16'hFFFF;
rommem[9041] <= 16'hFFFF;
rommem[9042] <= 16'hFFFF;
rommem[9043] <= 16'hFFFF;
rommem[9044] <= 16'hFFFF;
rommem[9045] <= 16'hFFFF;
rommem[9046] <= 16'hFFFF;
rommem[9047] <= 16'hFFFF;
rommem[9048] <= 16'hFFFF;
rommem[9049] <= 16'hFFFF;
rommem[9050] <= 16'hFFFF;
rommem[9051] <= 16'hFFFF;
rommem[9052] <= 16'hFFFF;
rommem[9053] <= 16'hFFFF;
rommem[9054] <= 16'hFFFF;
rommem[9055] <= 16'hFFFF;
rommem[9056] <= 16'hFFFF;
rommem[9057] <= 16'hFFFF;
rommem[9058] <= 16'hFFFF;
rommem[9059] <= 16'hFFFF;
rommem[9060] <= 16'hFFFF;
rommem[9061] <= 16'hFFFF;
rommem[9062] <= 16'hFFFF;
rommem[9063] <= 16'hFFFF;
rommem[9064] <= 16'hFFFF;
rommem[9065] <= 16'hFFFF;
rommem[9066] <= 16'hFFFF;
rommem[9067] <= 16'hFFFF;
rommem[9068] <= 16'hFFFF;
rommem[9069] <= 16'hFFFF;
rommem[9070] <= 16'hFFFF;
rommem[9071] <= 16'hFFFF;
rommem[9072] <= 16'hFFFF;
rommem[9073] <= 16'hFFFF;
rommem[9074] <= 16'hFFFF;
rommem[9075] <= 16'hFFFF;
rommem[9076] <= 16'hFFFF;
rommem[9077] <= 16'hFFFF;
rommem[9078] <= 16'hFFFF;
rommem[9079] <= 16'hFFFF;
rommem[9080] <= 16'hFFFF;
rommem[9081] <= 16'hFFFF;
rommem[9082] <= 16'hFFFF;
rommem[9083] <= 16'hFFFF;
rommem[9084] <= 16'hFFFF;
rommem[9085] <= 16'hFFFF;
rommem[9086] <= 16'hFFFF;
rommem[9087] <= 16'hFFFF;
rommem[9088] <= 16'hFFFF;
rommem[9089] <= 16'hFFFF;
rommem[9090] <= 16'hFFFF;
rommem[9091] <= 16'hFFFF;
rommem[9092] <= 16'hFFFF;
rommem[9093] <= 16'hFFFF;
rommem[9094] <= 16'hFFFF;
rommem[9095] <= 16'hFFFF;
rommem[9096] <= 16'hFFFF;
rommem[9097] <= 16'hFFFF;
rommem[9098] <= 16'hFFFF;
rommem[9099] <= 16'hFFFF;
rommem[9100] <= 16'hFFFF;
rommem[9101] <= 16'hFFFF;
rommem[9102] <= 16'hFFFF;
rommem[9103] <= 16'hFFFF;
rommem[9104] <= 16'hFFFF;
rommem[9105] <= 16'hFFFF;
rommem[9106] <= 16'hFFFF;
rommem[9107] <= 16'hFFFF;
rommem[9108] <= 16'hFFFF;
rommem[9109] <= 16'hFFFF;
rommem[9110] <= 16'hFFFF;
rommem[9111] <= 16'hFFFF;
rommem[9112] <= 16'hFFFF;
rommem[9113] <= 16'hFFFF;
rommem[9114] <= 16'hFFFF;
rommem[9115] <= 16'hFFFF;
rommem[9116] <= 16'hFFFF;
rommem[9117] <= 16'hFFFF;
rommem[9118] <= 16'hFFFF;
rommem[9119] <= 16'hFFFF;
rommem[9120] <= 16'hFFFF;
rommem[9121] <= 16'hFFFF;
rommem[9122] <= 16'hFFFF;
rommem[9123] <= 16'hFFFF;
rommem[9124] <= 16'hFFFF;
rommem[9125] <= 16'hFFFF;
rommem[9126] <= 16'hFFFF;
rommem[9127] <= 16'hFFFF;
rommem[9128] <= 16'hFFFF;
rommem[9129] <= 16'hFFFF;
rommem[9130] <= 16'hFFFF;
rommem[9131] <= 16'hFFFF;
rommem[9132] <= 16'hFFFF;
rommem[9133] <= 16'hFFFF;
rommem[9134] <= 16'hFFFF;
rommem[9135] <= 16'hFFFF;
rommem[9136] <= 16'hFFFF;
rommem[9137] <= 16'hFFFF;
rommem[9138] <= 16'hFFFF;
rommem[9139] <= 16'hFFFF;
rommem[9140] <= 16'hFFFF;
rommem[9141] <= 16'hFFFF;
rommem[9142] <= 16'hFFFF;
rommem[9143] <= 16'hFFFF;
rommem[9144] <= 16'hFFFF;
rommem[9145] <= 16'hFFFF;
rommem[9146] <= 16'hFFFF;
rommem[9147] <= 16'hFFFF;
rommem[9148] <= 16'hFFFF;
rommem[9149] <= 16'hFFFF;
rommem[9150] <= 16'hFFFF;
rommem[9151] <= 16'hFFFF;
rommem[9152] <= 16'hFFFF;
rommem[9153] <= 16'hFFFF;
rommem[9154] <= 16'hFFFF;
rommem[9155] <= 16'hFFFF;
rommem[9156] <= 16'hFFFF;
rommem[9157] <= 16'hFFFF;
rommem[9158] <= 16'hFFFF;
rommem[9159] <= 16'hFFFF;
rommem[9160] <= 16'hFFFF;
rommem[9161] <= 16'hFFFF;
rommem[9162] <= 16'hFFFF;
rommem[9163] <= 16'hFFFF;
rommem[9164] <= 16'hFFFF;
rommem[9165] <= 16'hFFFF;
rommem[9166] <= 16'hFFFF;
rommem[9167] <= 16'hFFFF;
rommem[9168] <= 16'hFFFF;
rommem[9169] <= 16'hFFFF;
rommem[9170] <= 16'hFFFF;
rommem[9171] <= 16'hFFFF;
rommem[9172] <= 16'hFFFF;
rommem[9173] <= 16'hFFFF;
rommem[9174] <= 16'hFFFF;
rommem[9175] <= 16'hFFFF;
rommem[9176] <= 16'hFFFF;
rommem[9177] <= 16'hFFFF;
rommem[9178] <= 16'hFFFF;
rommem[9179] <= 16'hFFFF;
rommem[9180] <= 16'hFFFF;
rommem[9181] <= 16'hFFFF;
rommem[9182] <= 16'hFFFF;
rommem[9183] <= 16'hFFFF;
rommem[9184] <= 16'hFFFF;
rommem[9185] <= 16'hFFFF;
rommem[9186] <= 16'hFFFF;
rommem[9187] <= 16'hFFFF;
rommem[9188] <= 16'hFFFF;
rommem[9189] <= 16'hFFFF;
rommem[9190] <= 16'hFFFF;
rommem[9191] <= 16'hFFFF;
rommem[9192] <= 16'hFFFF;
rommem[9193] <= 16'hFFFF;
rommem[9194] <= 16'hFFFF;
rommem[9195] <= 16'hFFFF;
rommem[9196] <= 16'hFFFF;
rommem[9197] <= 16'hFFFF;
rommem[9198] <= 16'hFFFF;
rommem[9199] <= 16'hFFFF;
rommem[9200] <= 16'hFFFF;
rommem[9201] <= 16'hFFFF;
rommem[9202] <= 16'hFFFF;
rommem[9203] <= 16'hFFFF;
rommem[9204] <= 16'hFFFF;
rommem[9205] <= 16'hFFFF;
rommem[9206] <= 16'hFFFF;
rommem[9207] <= 16'hFFFF;
rommem[9208] <= 16'hFFFF;
rommem[9209] <= 16'hFFFF;
rommem[9210] <= 16'hFFFF;
rommem[9211] <= 16'hFFFF;
rommem[9212] <= 16'hFFFF;
rommem[9213] <= 16'hFFFF;
rommem[9214] <= 16'hFFFF;
rommem[9215] <= 16'hFFFF;
rommem[9216] <= 16'hFFFF;
rommem[9217] <= 16'hFFFF;
rommem[9218] <= 16'hFFFF;
rommem[9219] <= 16'hFFFF;
rommem[9220] <= 16'hFFFF;
rommem[9221] <= 16'hFFFF;
rommem[9222] <= 16'hFFFF;
rommem[9223] <= 16'hFFFF;
rommem[9224] <= 16'hFFFF;
rommem[9225] <= 16'hFFFF;
rommem[9226] <= 16'hFFFF;
rommem[9227] <= 16'hFFFF;
rommem[9228] <= 16'hFFFF;
rommem[9229] <= 16'hFFFF;
rommem[9230] <= 16'hFFFF;
rommem[9231] <= 16'hFFFF;
rommem[9232] <= 16'hFFFF;
rommem[9233] <= 16'hFFFF;
rommem[9234] <= 16'hFFFF;
rommem[9235] <= 16'hFFFF;
rommem[9236] <= 16'hFFFF;
rommem[9237] <= 16'hFFFF;
rommem[9238] <= 16'hFFFF;
rommem[9239] <= 16'hFFFF;
rommem[9240] <= 16'hFFFF;
rommem[9241] <= 16'hFFFF;
rommem[9242] <= 16'hFFFF;
rommem[9243] <= 16'hFFFF;
rommem[9244] <= 16'hFFFF;
rommem[9245] <= 16'hFFFF;
rommem[9246] <= 16'hFFFF;
rommem[9247] <= 16'hFFFF;
rommem[9248] <= 16'hFFFF;
rommem[9249] <= 16'hFFFF;
rommem[9250] <= 16'hFFFF;
rommem[9251] <= 16'hFFFF;
rommem[9252] <= 16'hFFFF;
rommem[9253] <= 16'hFFFF;
rommem[9254] <= 16'hFFFF;
rommem[9255] <= 16'hFFFF;
rommem[9256] <= 16'hFFFF;
rommem[9257] <= 16'hFFFF;
rommem[9258] <= 16'hFFFF;
rommem[9259] <= 16'hFFFF;
rommem[9260] <= 16'hFFFF;
rommem[9261] <= 16'hFFFF;
rommem[9262] <= 16'hFFFF;
rommem[9263] <= 16'hFFFF;
rommem[9264] <= 16'hFFFF;
rommem[9265] <= 16'hFFFF;
rommem[9266] <= 16'hFFFF;
rommem[9267] <= 16'hFFFF;
rommem[9268] <= 16'hFFFF;
rommem[9269] <= 16'hFFFF;
rommem[9270] <= 16'hFFFF;
rommem[9271] <= 16'hFFFF;
rommem[9272] <= 16'hFFFF;
rommem[9273] <= 16'hFFFF;
rommem[9274] <= 16'hFFFF;
rommem[9275] <= 16'hFFFF;
rommem[9276] <= 16'hFFFF;
rommem[9277] <= 16'hFFFF;
rommem[9278] <= 16'hFFFF;
rommem[9279] <= 16'hFFFF;
rommem[9280] <= 16'hFFFF;
rommem[9281] <= 16'hFFFF;
rommem[9282] <= 16'hFFFF;
rommem[9283] <= 16'hFFFF;
rommem[9284] <= 16'hFFFF;
rommem[9285] <= 16'hFFFF;
rommem[9286] <= 16'hFFFF;
rommem[9287] <= 16'hFFFF;
rommem[9288] <= 16'hFFFF;
rommem[9289] <= 16'hFFFF;
rommem[9290] <= 16'hFFFF;
rommem[9291] <= 16'hFFFF;
rommem[9292] <= 16'hFFFF;
rommem[9293] <= 16'hFFFF;
rommem[9294] <= 16'hFFFF;
rommem[9295] <= 16'hFFFF;
rommem[9296] <= 16'hFFFF;
rommem[9297] <= 16'hFFFF;
rommem[9298] <= 16'hFFFF;
rommem[9299] <= 16'hFFFF;
rommem[9300] <= 16'hFFFF;
rommem[9301] <= 16'hFFFF;
rommem[9302] <= 16'hFFFF;
rommem[9303] <= 16'hFFFF;
rommem[9304] <= 16'hFFFF;
rommem[9305] <= 16'hFFFF;
rommem[9306] <= 16'hFFFF;
rommem[9307] <= 16'hFFFF;
rommem[9308] <= 16'hFFFF;
rommem[9309] <= 16'hFFFF;
rommem[9310] <= 16'hFFFF;
rommem[9311] <= 16'hFFFF;
rommem[9312] <= 16'hFFFF;
rommem[9313] <= 16'hFFFF;
rommem[9314] <= 16'hFFFF;
rommem[9315] <= 16'hFFFF;
rommem[9316] <= 16'hFFFF;
rommem[9317] <= 16'hFFFF;
rommem[9318] <= 16'hFFFF;
rommem[9319] <= 16'hFFFF;
rommem[9320] <= 16'hFFFF;
rommem[9321] <= 16'hFFFF;
rommem[9322] <= 16'hFFFF;
rommem[9323] <= 16'hFFFF;
rommem[9324] <= 16'hFFFF;
rommem[9325] <= 16'hFFFF;
rommem[9326] <= 16'hFFFF;
rommem[9327] <= 16'hFFFF;
rommem[9328] <= 16'hFFFF;
rommem[9329] <= 16'hFFFF;
rommem[9330] <= 16'hFFFF;
rommem[9331] <= 16'hFFFF;
rommem[9332] <= 16'hFFFF;
rommem[9333] <= 16'hFFFF;
rommem[9334] <= 16'hFFFF;
rommem[9335] <= 16'hFFFF;
rommem[9336] <= 16'hFFFF;
rommem[9337] <= 16'hFFFF;
rommem[9338] <= 16'hFFFF;
rommem[9339] <= 16'hFFFF;
rommem[9340] <= 16'hFFFF;
rommem[9341] <= 16'hFFFF;
rommem[9342] <= 16'hFFFF;
rommem[9343] <= 16'hFFFF;
rommem[9344] <= 16'hFFFF;
rommem[9345] <= 16'hFFFF;
rommem[9346] <= 16'hFFFF;
rommem[9347] <= 16'hFFFF;
rommem[9348] <= 16'hFFFF;
rommem[9349] <= 16'hFFFF;
rommem[9350] <= 16'hFFFF;
rommem[9351] <= 16'hFFFF;
rommem[9352] <= 16'hFFFF;
rommem[9353] <= 16'hFFFF;
rommem[9354] <= 16'hFFFF;
rommem[9355] <= 16'hFFFF;
rommem[9356] <= 16'hFFFF;
rommem[9357] <= 16'hFFFF;
rommem[9358] <= 16'hFFFF;
rommem[9359] <= 16'hFFFF;
rommem[9360] <= 16'hFFFF;
rommem[9361] <= 16'hFFFF;
rommem[9362] <= 16'hFFFF;
rommem[9363] <= 16'hFFFF;
rommem[9364] <= 16'hFFFF;
rommem[9365] <= 16'hFFFF;
rommem[9366] <= 16'hFFFF;
rommem[9367] <= 16'hFFFF;
rommem[9368] <= 16'hFFFF;
rommem[9369] <= 16'hFFFF;
rommem[9370] <= 16'hFFFF;
rommem[9371] <= 16'hFFFF;
rommem[9372] <= 16'hFFFF;
rommem[9373] <= 16'hFFFF;
rommem[9374] <= 16'hFFFF;
rommem[9375] <= 16'hFFFF;
rommem[9376] <= 16'hFFFF;
rommem[9377] <= 16'hFFFF;
rommem[9378] <= 16'hFFFF;
rommem[9379] <= 16'hFFFF;
rommem[9380] <= 16'hFFFF;
rommem[9381] <= 16'hFFFF;
rommem[9382] <= 16'hFFFF;
rommem[9383] <= 16'hFFFF;
rommem[9384] <= 16'hFFFF;
rommem[9385] <= 16'hFFFF;
rommem[9386] <= 16'hFFFF;
rommem[9387] <= 16'hFFFF;
rommem[9388] <= 16'hFFFF;
rommem[9389] <= 16'hFFFF;
rommem[9390] <= 16'hFFFF;
rommem[9391] <= 16'hFFFF;
rommem[9392] <= 16'hFFFF;
rommem[9393] <= 16'hFFFF;
rommem[9394] <= 16'hFFFF;
rommem[9395] <= 16'hFFFF;
rommem[9396] <= 16'hFFFF;
rommem[9397] <= 16'hFFFF;
rommem[9398] <= 16'hFFFF;
rommem[9399] <= 16'hFFFF;
rommem[9400] <= 16'hFFFF;
rommem[9401] <= 16'hFFFF;
rommem[9402] <= 16'hFFFF;
rommem[9403] <= 16'hFFFF;
rommem[9404] <= 16'hFFFF;
rommem[9405] <= 16'hFFFF;
rommem[9406] <= 16'hFFFF;
rommem[9407] <= 16'hFFFF;
rommem[9408] <= 16'hFFFF;
rommem[9409] <= 16'hFFFF;
rommem[9410] <= 16'hFFFF;
rommem[9411] <= 16'hFFFF;
rommem[9412] <= 16'hFFFF;
rommem[9413] <= 16'hFFFF;
rommem[9414] <= 16'hFFFF;
rommem[9415] <= 16'hFFFF;
rommem[9416] <= 16'hFFFF;
rommem[9417] <= 16'hFFFF;
rommem[9418] <= 16'hFFFF;
rommem[9419] <= 16'hFFFF;
rommem[9420] <= 16'hFFFF;
rommem[9421] <= 16'hFFFF;
rommem[9422] <= 16'hFFFF;
rommem[9423] <= 16'hFFFF;
rommem[9424] <= 16'hFFFF;
rommem[9425] <= 16'hFFFF;
rommem[9426] <= 16'hFFFF;
rommem[9427] <= 16'hFFFF;
rommem[9428] <= 16'hFFFF;
rommem[9429] <= 16'hFFFF;
rommem[9430] <= 16'hFFFF;
rommem[9431] <= 16'hFFFF;
rommem[9432] <= 16'hFFFF;
rommem[9433] <= 16'hFFFF;
rommem[9434] <= 16'hFFFF;
rommem[9435] <= 16'hFFFF;
rommem[9436] <= 16'hFFFF;
rommem[9437] <= 16'hFFFF;
rommem[9438] <= 16'hFFFF;
rommem[9439] <= 16'hFFFF;
rommem[9440] <= 16'hFFFF;
rommem[9441] <= 16'hFFFF;
rommem[9442] <= 16'hFFFF;
rommem[9443] <= 16'hFFFF;
rommem[9444] <= 16'hFFFF;
rommem[9445] <= 16'hFFFF;
rommem[9446] <= 16'hFFFF;
rommem[9447] <= 16'hFFFF;
rommem[9448] <= 16'hFFFF;
rommem[9449] <= 16'hFFFF;
rommem[9450] <= 16'hFFFF;
rommem[9451] <= 16'hFFFF;
rommem[9452] <= 16'hFFFF;
rommem[9453] <= 16'hFFFF;
rommem[9454] <= 16'hFFFF;
rommem[9455] <= 16'hFFFF;
rommem[9456] <= 16'hFFFF;
rommem[9457] <= 16'hFFFF;
rommem[9458] <= 16'hFFFF;
rommem[9459] <= 16'hFFFF;
rommem[9460] <= 16'hFFFF;
rommem[9461] <= 16'hFFFF;
rommem[9462] <= 16'hFFFF;
rommem[9463] <= 16'hFFFF;
rommem[9464] <= 16'hFFFF;
rommem[9465] <= 16'hFFFF;
rommem[9466] <= 16'hFFFF;
rommem[9467] <= 16'hFFFF;
rommem[9468] <= 16'hFFFF;
rommem[9469] <= 16'hFFFF;
rommem[9470] <= 16'hFFFF;
rommem[9471] <= 16'hFFFF;
rommem[9472] <= 16'hFFFF;
rommem[9473] <= 16'hFFFF;
rommem[9474] <= 16'hFFFF;
rommem[9475] <= 16'hFFFF;
rommem[9476] <= 16'hFFFF;
rommem[9477] <= 16'hFFFF;
rommem[9478] <= 16'hFFFF;
rommem[9479] <= 16'hFFFF;
rommem[9480] <= 16'hFFFF;
rommem[9481] <= 16'hFFFF;
rommem[9482] <= 16'hFFFF;
rommem[9483] <= 16'hFFFF;
rommem[9484] <= 16'hFFFF;
rommem[9485] <= 16'hFFFF;
rommem[9486] <= 16'hFFFF;
rommem[9487] <= 16'hFFFF;
rommem[9488] <= 16'hFFFF;
rommem[9489] <= 16'hFFFF;
rommem[9490] <= 16'hFFFF;
rommem[9491] <= 16'hFFFF;
rommem[9492] <= 16'hFFFF;
rommem[9493] <= 16'hFFFF;
rommem[9494] <= 16'hFFFF;
rommem[9495] <= 16'hFFFF;
rommem[9496] <= 16'hFFFF;
rommem[9497] <= 16'hFFFF;
rommem[9498] <= 16'hFFFF;
rommem[9499] <= 16'hFFFF;
rommem[9500] <= 16'hFFFF;
rommem[9501] <= 16'hFFFF;
rommem[9502] <= 16'hFFFF;
rommem[9503] <= 16'hFFFF;
rommem[9504] <= 16'hFFFF;
rommem[9505] <= 16'hFFFF;
rommem[9506] <= 16'hFFFF;
rommem[9507] <= 16'hFFFF;
rommem[9508] <= 16'hFFFF;
rommem[9509] <= 16'hFFFF;
rommem[9510] <= 16'hFFFF;
rommem[9511] <= 16'hFFFF;
rommem[9512] <= 16'hFFFF;
rommem[9513] <= 16'hFFFF;
rommem[9514] <= 16'hFFFF;
rommem[9515] <= 16'hFFFF;
rommem[9516] <= 16'hFFFF;
rommem[9517] <= 16'hFFFF;
rommem[9518] <= 16'hFFFF;
rommem[9519] <= 16'hFFFF;
rommem[9520] <= 16'hFFFF;
rommem[9521] <= 16'hFFFF;
rommem[9522] <= 16'hFFFF;
rommem[9523] <= 16'hFFFF;
rommem[9524] <= 16'hFFFF;
rommem[9525] <= 16'hFFFF;
rommem[9526] <= 16'hFFFF;
rommem[9527] <= 16'hFFFF;
rommem[9528] <= 16'hFFFF;
rommem[9529] <= 16'hFFFF;
rommem[9530] <= 16'hFFFF;
rommem[9531] <= 16'hFFFF;
rommem[9532] <= 16'hFFFF;
rommem[9533] <= 16'hFFFF;
rommem[9534] <= 16'hFFFF;
rommem[9535] <= 16'hFFFF;
rommem[9536] <= 16'hFFFF;
rommem[9537] <= 16'hFFFF;
rommem[9538] <= 16'hFFFF;
rommem[9539] <= 16'hFFFF;
rommem[9540] <= 16'hFFFF;
rommem[9541] <= 16'hFFFF;
rommem[9542] <= 16'hFFFF;
rommem[9543] <= 16'hFFFF;
rommem[9544] <= 16'hFFFF;
rommem[9545] <= 16'hFFFF;
rommem[9546] <= 16'hFFFF;
rommem[9547] <= 16'hFFFF;
rommem[9548] <= 16'hFFFF;
rommem[9549] <= 16'hFFFF;
rommem[9550] <= 16'hFFFF;
rommem[9551] <= 16'hFFFF;
rommem[9552] <= 16'hFFFF;
rommem[9553] <= 16'hFFFF;
rommem[9554] <= 16'hFFFF;
rommem[9555] <= 16'hFFFF;
rommem[9556] <= 16'hFFFF;
rommem[9557] <= 16'hFFFF;
rommem[9558] <= 16'hFFFF;
rommem[9559] <= 16'hFFFF;
rommem[9560] <= 16'hFFFF;
rommem[9561] <= 16'hFFFF;
rommem[9562] <= 16'hFFFF;
rommem[9563] <= 16'hFFFF;
rommem[9564] <= 16'hFFFF;
rommem[9565] <= 16'hFFFF;
rommem[9566] <= 16'hFFFF;
rommem[9567] <= 16'hFFFF;
rommem[9568] <= 16'hFFFF;
rommem[9569] <= 16'hFFFF;
rommem[9570] <= 16'hFFFF;
rommem[9571] <= 16'hFFFF;
rommem[9572] <= 16'hFFFF;
rommem[9573] <= 16'hFFFF;
rommem[9574] <= 16'hFFFF;
rommem[9575] <= 16'hFFFF;
rommem[9576] <= 16'hFFFF;
rommem[9577] <= 16'hFFFF;
rommem[9578] <= 16'hFFFF;
rommem[9579] <= 16'hFFFF;
rommem[9580] <= 16'hFFFF;
rommem[9581] <= 16'hFFFF;
rommem[9582] <= 16'hFFFF;
rommem[9583] <= 16'hFFFF;
rommem[9584] <= 16'hFFFF;
rommem[9585] <= 16'hFFFF;
rommem[9586] <= 16'hFFFF;
rommem[9587] <= 16'hFFFF;
rommem[9588] <= 16'hFFFF;
rommem[9589] <= 16'hFFFF;
rommem[9590] <= 16'hFFFF;
rommem[9591] <= 16'hFFFF;
rommem[9592] <= 16'hFFFF;
rommem[9593] <= 16'hFFFF;
rommem[9594] <= 16'hFFFF;
rommem[9595] <= 16'hFFFF;
rommem[9596] <= 16'hFFFF;
rommem[9597] <= 16'hFFFF;
rommem[9598] <= 16'hFFFF;
rommem[9599] <= 16'hFFFF;
rommem[9600] <= 16'hFFFF;
rommem[9601] <= 16'hFFFF;
rommem[9602] <= 16'hFFFF;
rommem[9603] <= 16'hFFFF;
rommem[9604] <= 16'hFFFF;
rommem[9605] <= 16'hFFFF;
rommem[9606] <= 16'hFFFF;
rommem[9607] <= 16'hFFFF;
rommem[9608] <= 16'hFFFF;
rommem[9609] <= 16'hFFFF;
rommem[9610] <= 16'hFFFF;
rommem[9611] <= 16'hFFFF;
rommem[9612] <= 16'hFFFF;
rommem[9613] <= 16'hFFFF;
rommem[9614] <= 16'hFFFF;
rommem[9615] <= 16'hFFFF;
rommem[9616] <= 16'hFFFF;
rommem[9617] <= 16'hFFFF;
rommem[9618] <= 16'hFFFF;
rommem[9619] <= 16'hFFFF;
rommem[9620] <= 16'hFFFF;
rommem[9621] <= 16'hFFFF;
rommem[9622] <= 16'hFFFF;
rommem[9623] <= 16'hFFFF;
rommem[9624] <= 16'hFFFF;
rommem[9625] <= 16'hFFFF;
rommem[9626] <= 16'hFFFF;
rommem[9627] <= 16'hFFFF;
rommem[9628] <= 16'hFFFF;
rommem[9629] <= 16'hFFFF;
rommem[9630] <= 16'hFFFF;
rommem[9631] <= 16'hFFFF;
rommem[9632] <= 16'hFFFF;
rommem[9633] <= 16'hFFFF;
rommem[9634] <= 16'hFFFF;
rommem[9635] <= 16'hFFFF;
rommem[9636] <= 16'hFFFF;
rommem[9637] <= 16'hFFFF;
rommem[9638] <= 16'hFFFF;
rommem[9639] <= 16'hFFFF;
rommem[9640] <= 16'hFFFF;
rommem[9641] <= 16'hFFFF;
rommem[9642] <= 16'hFFFF;
rommem[9643] <= 16'hFFFF;
rommem[9644] <= 16'hFFFF;
rommem[9645] <= 16'hFFFF;
rommem[9646] <= 16'hFFFF;
rommem[9647] <= 16'hFFFF;
rommem[9648] <= 16'hFFFF;
rommem[9649] <= 16'hFFFF;
rommem[9650] <= 16'hFFFF;
rommem[9651] <= 16'hFFFF;
rommem[9652] <= 16'hFFFF;
rommem[9653] <= 16'hFFFF;
rommem[9654] <= 16'hFFFF;
rommem[9655] <= 16'hFFFF;
rommem[9656] <= 16'hFFFF;
rommem[9657] <= 16'hFFFF;
rommem[9658] <= 16'hFFFF;
rommem[9659] <= 16'hFFFF;
rommem[9660] <= 16'hFFFF;
rommem[9661] <= 16'hFFFF;
rommem[9662] <= 16'hFFFF;
rommem[9663] <= 16'hFFFF;
rommem[9664] <= 16'hFFFF;
rommem[9665] <= 16'hFFFF;
rommem[9666] <= 16'hFFFF;
rommem[9667] <= 16'hFFFF;
rommem[9668] <= 16'hFFFF;
rommem[9669] <= 16'hFFFF;
rommem[9670] <= 16'hFFFF;
rommem[9671] <= 16'hFFFF;
rommem[9672] <= 16'hFFFF;
rommem[9673] <= 16'hFFFF;
rommem[9674] <= 16'hFFFF;
rommem[9675] <= 16'hFFFF;
rommem[9676] <= 16'hFFFF;
rommem[9677] <= 16'hFFFF;
rommem[9678] <= 16'hFFFF;
rommem[9679] <= 16'hFFFF;
rommem[9680] <= 16'hFFFF;
rommem[9681] <= 16'hFFFF;
rommem[9682] <= 16'hFFFF;
rommem[9683] <= 16'hFFFF;
rommem[9684] <= 16'hFFFF;
rommem[9685] <= 16'hFFFF;
rommem[9686] <= 16'hFFFF;
rommem[9687] <= 16'hFFFF;
rommem[9688] <= 16'hFFFF;
rommem[9689] <= 16'hFFFF;
rommem[9690] <= 16'hFFFF;
rommem[9691] <= 16'hFFFF;
rommem[9692] <= 16'hFFFF;
rommem[9693] <= 16'hFFFF;
rommem[9694] <= 16'hFFFF;
rommem[9695] <= 16'hFFFF;
rommem[9696] <= 16'hFFFF;
rommem[9697] <= 16'hFFFF;
rommem[9698] <= 16'hFFFF;
rommem[9699] <= 16'hFFFF;
rommem[9700] <= 16'hFFFF;
rommem[9701] <= 16'hFFFF;
rommem[9702] <= 16'hFFFF;
rommem[9703] <= 16'hFFFF;
rommem[9704] <= 16'hFFFF;
rommem[9705] <= 16'hFFFF;
rommem[9706] <= 16'hFFFF;
rommem[9707] <= 16'hFFFF;
rommem[9708] <= 16'hFFFF;
rommem[9709] <= 16'hFFFF;
rommem[9710] <= 16'hFFFF;
rommem[9711] <= 16'hFFFF;
rommem[9712] <= 16'hFFFF;
rommem[9713] <= 16'hFFFF;
rommem[9714] <= 16'hFFFF;
rommem[9715] <= 16'hFFFF;
rommem[9716] <= 16'hFFFF;
rommem[9717] <= 16'hFFFF;
rommem[9718] <= 16'hFFFF;
rommem[9719] <= 16'hFFFF;
rommem[9720] <= 16'hFFFF;
rommem[9721] <= 16'hFFFF;
rommem[9722] <= 16'hFFFF;
rommem[9723] <= 16'hFFFF;
rommem[9724] <= 16'hFFFF;
rommem[9725] <= 16'hFFFF;
rommem[9726] <= 16'hFFFF;
rommem[9727] <= 16'hFFFF;
rommem[9728] <= 16'hFFFF;
rommem[9729] <= 16'hFFFF;
rommem[9730] <= 16'hFFFF;
rommem[9731] <= 16'hFFFF;
rommem[9732] <= 16'hFFFF;
rommem[9733] <= 16'hFFFF;
rommem[9734] <= 16'hFFFF;
rommem[9735] <= 16'hFFFF;
rommem[9736] <= 16'hFFFF;
rommem[9737] <= 16'hFFFF;
rommem[9738] <= 16'hFFFF;
rommem[9739] <= 16'hFFFF;
rommem[9740] <= 16'hFFFF;
rommem[9741] <= 16'hFFFF;
rommem[9742] <= 16'hFFFF;
rommem[9743] <= 16'hFFFF;
rommem[9744] <= 16'hFFFF;
rommem[9745] <= 16'hFFFF;
rommem[9746] <= 16'hFFFF;
rommem[9747] <= 16'hFFFF;
rommem[9748] <= 16'hFFFF;
rommem[9749] <= 16'hFFFF;
rommem[9750] <= 16'hFFFF;
rommem[9751] <= 16'hFFFF;
rommem[9752] <= 16'hFFFF;
rommem[9753] <= 16'hFFFF;
rommem[9754] <= 16'hFFFF;
rommem[9755] <= 16'hFFFF;
rommem[9756] <= 16'hFFFF;
rommem[9757] <= 16'hFFFF;
rommem[9758] <= 16'hFFFF;
rommem[9759] <= 16'hFFFF;
rommem[9760] <= 16'hFFFF;
rommem[9761] <= 16'hFFFF;
rommem[9762] <= 16'hFFFF;
rommem[9763] <= 16'hFFFF;
rommem[9764] <= 16'hFFFF;
rommem[9765] <= 16'hFFFF;
rommem[9766] <= 16'hFFFF;
rommem[9767] <= 16'hFFFF;
rommem[9768] <= 16'hFFFF;
rommem[9769] <= 16'hFFFF;
rommem[9770] <= 16'hFFFF;
rommem[9771] <= 16'hFFFF;
rommem[9772] <= 16'hFFFF;
rommem[9773] <= 16'hFFFF;
rommem[9774] <= 16'hFFFF;
rommem[9775] <= 16'hFFFF;
rommem[9776] <= 16'hFFFF;
rommem[9777] <= 16'hFFFF;
rommem[9778] <= 16'hFFFF;
rommem[9779] <= 16'hFFFF;
rommem[9780] <= 16'hFFFF;
rommem[9781] <= 16'hFFFF;
rommem[9782] <= 16'hFFFF;
rommem[9783] <= 16'hFFFF;
rommem[9784] <= 16'hFFFF;
rommem[9785] <= 16'hFFFF;
rommem[9786] <= 16'hFFFF;
rommem[9787] <= 16'hFFFF;
rommem[9788] <= 16'hFFFF;
rommem[9789] <= 16'hFFFF;
rommem[9790] <= 16'hFFFF;
rommem[9791] <= 16'hFFFF;
rommem[9792] <= 16'hFFFF;
rommem[9793] <= 16'hFFFF;
rommem[9794] <= 16'hFFFF;
rommem[9795] <= 16'hFFFF;
rommem[9796] <= 16'hFFFF;
rommem[9797] <= 16'hFFFF;
rommem[9798] <= 16'hFFFF;
rommem[9799] <= 16'hFFFF;
rommem[9800] <= 16'hFFFF;
rommem[9801] <= 16'hFFFF;
rommem[9802] <= 16'hFFFF;
rommem[9803] <= 16'hFFFF;
rommem[9804] <= 16'hFFFF;
rommem[9805] <= 16'hFFFF;
rommem[9806] <= 16'hFFFF;
rommem[9807] <= 16'hFFFF;
rommem[9808] <= 16'hFFFF;
rommem[9809] <= 16'hFFFF;
rommem[9810] <= 16'hFFFF;
rommem[9811] <= 16'hFFFF;
rommem[9812] <= 16'hFFFF;
rommem[9813] <= 16'hFFFF;
rommem[9814] <= 16'hFFFF;
rommem[9815] <= 16'hFFFF;
rommem[9816] <= 16'hFFFF;
rommem[9817] <= 16'hFFFF;
rommem[9818] <= 16'hFFFF;
rommem[9819] <= 16'hFFFF;
rommem[9820] <= 16'hFFFF;
rommem[9821] <= 16'hFFFF;
rommem[9822] <= 16'hFFFF;
rommem[9823] <= 16'hFFFF;
rommem[9824] <= 16'hFFFF;
rommem[9825] <= 16'hFFFF;
rommem[9826] <= 16'hFFFF;
rommem[9827] <= 16'hFFFF;
rommem[9828] <= 16'hFFFF;
rommem[9829] <= 16'hFFFF;
rommem[9830] <= 16'hFFFF;
rommem[9831] <= 16'hFFFF;
rommem[9832] <= 16'hFFFF;
rommem[9833] <= 16'hFFFF;
rommem[9834] <= 16'hFFFF;
rommem[9835] <= 16'hFFFF;
rommem[9836] <= 16'hFFFF;
rommem[9837] <= 16'hFFFF;
rommem[9838] <= 16'hFFFF;
rommem[9839] <= 16'hFFFF;
rommem[9840] <= 16'hFFFF;
rommem[9841] <= 16'hFFFF;
rommem[9842] <= 16'hFFFF;
rommem[9843] <= 16'hFFFF;
rommem[9844] <= 16'hFFFF;
rommem[9845] <= 16'hFFFF;
rommem[9846] <= 16'hFFFF;
rommem[9847] <= 16'hFFFF;
rommem[9848] <= 16'hFFFF;
rommem[9849] <= 16'hFFFF;
rommem[9850] <= 16'hFFFF;
rommem[9851] <= 16'hFFFF;
rommem[9852] <= 16'hFFFF;
rommem[9853] <= 16'hFFFF;
rommem[9854] <= 16'hFFFF;
rommem[9855] <= 16'hFFFF;
rommem[9856] <= 16'hFFFF;
rommem[9857] <= 16'hFFFF;
rommem[9858] <= 16'hFFFF;
rommem[9859] <= 16'hFFFF;
rommem[9860] <= 16'hFFFF;
rommem[9861] <= 16'hFFFF;
rommem[9862] <= 16'hFFFF;
rommem[9863] <= 16'hFFFF;
rommem[9864] <= 16'hFFFF;
rommem[9865] <= 16'hFFFF;
rommem[9866] <= 16'hFFFF;
rommem[9867] <= 16'hFFFF;
rommem[9868] <= 16'hFFFF;
rommem[9869] <= 16'hFFFF;
rommem[9870] <= 16'hFFFF;
rommem[9871] <= 16'hFFFF;
rommem[9872] <= 16'hFFFF;
rommem[9873] <= 16'hFFFF;
rommem[9874] <= 16'hFFFF;
rommem[9875] <= 16'hFFFF;
rommem[9876] <= 16'hFFFF;
rommem[9877] <= 16'hFFFF;
rommem[9878] <= 16'hFFFF;
rommem[9879] <= 16'hFFFF;
rommem[9880] <= 16'hFFFF;
rommem[9881] <= 16'hFFFF;
rommem[9882] <= 16'hFFFF;
rommem[9883] <= 16'hFFFF;
rommem[9884] <= 16'hFFFF;
rommem[9885] <= 16'hFFFF;
rommem[9886] <= 16'hFFFF;
rommem[9887] <= 16'hFFFF;
rommem[9888] <= 16'hFFFF;
rommem[9889] <= 16'hFFFF;
rommem[9890] <= 16'hFFFF;
rommem[9891] <= 16'hFFFF;
rommem[9892] <= 16'hFFFF;
rommem[9893] <= 16'hFFFF;
rommem[9894] <= 16'hFFFF;
rommem[9895] <= 16'hFFFF;
rommem[9896] <= 16'hFFFF;
rommem[9897] <= 16'hFFFF;
rommem[9898] <= 16'hFFFF;
rommem[9899] <= 16'hFFFF;
rommem[9900] <= 16'hFFFF;
rommem[9901] <= 16'hFFFF;
rommem[9902] <= 16'hFFFF;
rommem[9903] <= 16'hFFFF;
rommem[9904] <= 16'hFFFF;
rommem[9905] <= 16'hFFFF;
rommem[9906] <= 16'hFFFF;
rommem[9907] <= 16'hFFFF;
rommem[9908] <= 16'hFFFF;
rommem[9909] <= 16'hFFFF;
rommem[9910] <= 16'hFFFF;
rommem[9911] <= 16'hFFFF;
rommem[9912] <= 16'hFFFF;
rommem[9913] <= 16'hFFFF;
rommem[9914] <= 16'hFFFF;
rommem[9915] <= 16'hFFFF;
rommem[9916] <= 16'hFFFF;
rommem[9917] <= 16'hFFFF;
rommem[9918] <= 16'hFFFF;
rommem[9919] <= 16'hFFFF;
rommem[9920] <= 16'hFFFF;
rommem[9921] <= 16'hFFFF;
rommem[9922] <= 16'hFFFF;
rommem[9923] <= 16'hFFFF;
rommem[9924] <= 16'hFFFF;
rommem[9925] <= 16'hFFFF;
rommem[9926] <= 16'hFFFF;
rommem[9927] <= 16'hFFFF;
rommem[9928] <= 16'hFFFF;
rommem[9929] <= 16'hFFFF;
rommem[9930] <= 16'hFFFF;
rommem[9931] <= 16'hFFFF;
rommem[9932] <= 16'hFFFF;
rommem[9933] <= 16'hFFFF;
rommem[9934] <= 16'hFFFF;
rommem[9935] <= 16'hFFFF;
rommem[9936] <= 16'hFFFF;
rommem[9937] <= 16'hFFFF;
rommem[9938] <= 16'hFFFF;
rommem[9939] <= 16'hFFFF;
rommem[9940] <= 16'hFFFF;
rommem[9941] <= 16'hFFFF;
rommem[9942] <= 16'hFFFF;
rommem[9943] <= 16'hFFFF;
rommem[9944] <= 16'hFFFF;
rommem[9945] <= 16'hFFFF;
rommem[9946] <= 16'hFFFF;
rommem[9947] <= 16'hFFFF;
rommem[9948] <= 16'hFFFF;
rommem[9949] <= 16'hFFFF;
rommem[9950] <= 16'hFFFF;
rommem[9951] <= 16'hFFFF;
rommem[9952] <= 16'hFFFF;
rommem[9953] <= 16'hFFFF;
rommem[9954] <= 16'hFFFF;
rommem[9955] <= 16'hFFFF;
rommem[9956] <= 16'hFFFF;
rommem[9957] <= 16'hFFFF;
rommem[9958] <= 16'hFFFF;
rommem[9959] <= 16'hFFFF;
rommem[9960] <= 16'hFFFF;
rommem[9961] <= 16'hFFFF;
rommem[9962] <= 16'hFFFF;
rommem[9963] <= 16'hFFFF;
rommem[9964] <= 16'hFFFF;
rommem[9965] <= 16'hFFFF;
rommem[9966] <= 16'hFFFF;
rommem[9967] <= 16'hFFFF;
rommem[9968] <= 16'hFFFF;
rommem[9969] <= 16'hFFFF;
rommem[9970] <= 16'hFFFF;
rommem[9971] <= 16'hFFFF;
rommem[9972] <= 16'hFFFF;
rommem[9973] <= 16'hFFFF;
rommem[9974] <= 16'hFFFF;
rommem[9975] <= 16'hFFFF;
rommem[9976] <= 16'hFFFF;
rommem[9977] <= 16'hFFFF;
rommem[9978] <= 16'hFFFF;
rommem[9979] <= 16'hFFFF;
rommem[9980] <= 16'hFFFF;
rommem[9981] <= 16'hFFFF;
rommem[9982] <= 16'hFFFF;
rommem[9983] <= 16'hFFFF;
rommem[9984] <= 16'hFFFF;
rommem[9985] <= 16'hFFFF;
rommem[9986] <= 16'hFFFF;
rommem[9987] <= 16'hFFFF;
rommem[9988] <= 16'hFFFF;
rommem[9989] <= 16'hFFFF;
rommem[9990] <= 16'hFFFF;
rommem[9991] <= 16'hFFFF;
rommem[9992] <= 16'hFFFF;
rommem[9993] <= 16'hFFFF;
rommem[9994] <= 16'hFFFF;
rommem[9995] <= 16'hFFFF;
rommem[9996] <= 16'hFFFF;
rommem[9997] <= 16'hFFFF;
rommem[9998] <= 16'hFFFF;
rommem[9999] <= 16'hFFFF;
rommem[10000] <= 16'hFFFF;
rommem[10001] <= 16'hFFFF;
rommem[10002] <= 16'hFFFF;
rommem[10003] <= 16'hFFFF;
rommem[10004] <= 16'hFFFF;
rommem[10005] <= 16'hFFFF;
rommem[10006] <= 16'hFFFF;
rommem[10007] <= 16'hFFFF;
rommem[10008] <= 16'hFFFF;
rommem[10009] <= 16'hFFFF;
rommem[10010] <= 16'hFFFF;
rommem[10011] <= 16'hFFFF;
rommem[10012] <= 16'hFFFF;
rommem[10013] <= 16'hFFFF;
rommem[10014] <= 16'hFFFF;
rommem[10015] <= 16'hFFFF;
rommem[10016] <= 16'hFFFF;
rommem[10017] <= 16'hFFFF;
rommem[10018] <= 16'hFFFF;
rommem[10019] <= 16'hFFFF;
rommem[10020] <= 16'hFFFF;
rommem[10021] <= 16'hFFFF;
rommem[10022] <= 16'hFFFF;
rommem[10023] <= 16'hFFFF;
rommem[10024] <= 16'hFFFF;
rommem[10025] <= 16'hFFFF;
rommem[10026] <= 16'hFFFF;
rommem[10027] <= 16'hFFFF;
rommem[10028] <= 16'hFFFF;
rommem[10029] <= 16'hFFFF;
rommem[10030] <= 16'hFFFF;
rommem[10031] <= 16'hFFFF;
rommem[10032] <= 16'hFFFF;
rommem[10033] <= 16'hFFFF;
rommem[10034] <= 16'hFFFF;
rommem[10035] <= 16'hFFFF;
rommem[10036] <= 16'hFFFF;
rommem[10037] <= 16'hFFFF;
rommem[10038] <= 16'hFFFF;
rommem[10039] <= 16'hFFFF;
rommem[10040] <= 16'hFFFF;
rommem[10041] <= 16'hFFFF;
rommem[10042] <= 16'hFFFF;
rommem[10043] <= 16'hFFFF;
rommem[10044] <= 16'hFFFF;
rommem[10045] <= 16'hFFFF;
rommem[10046] <= 16'hFFFF;
rommem[10047] <= 16'hFFFF;
rommem[10048] <= 16'hFFFF;
rommem[10049] <= 16'hFFFF;
rommem[10050] <= 16'hFFFF;
rommem[10051] <= 16'hFFFF;
rommem[10052] <= 16'hFFFF;
rommem[10053] <= 16'hFFFF;
rommem[10054] <= 16'hFFFF;
rommem[10055] <= 16'hFFFF;
rommem[10056] <= 16'hFFFF;
rommem[10057] <= 16'hFFFF;
rommem[10058] <= 16'hFFFF;
rommem[10059] <= 16'hFFFF;
rommem[10060] <= 16'hFFFF;
rommem[10061] <= 16'hFFFF;
rommem[10062] <= 16'hFFFF;
rommem[10063] <= 16'hFFFF;
rommem[10064] <= 16'hFFFF;
rommem[10065] <= 16'hFFFF;
rommem[10066] <= 16'hFFFF;
rommem[10067] <= 16'hFFFF;
rommem[10068] <= 16'hFFFF;
rommem[10069] <= 16'hFFFF;
rommem[10070] <= 16'hFFFF;
rommem[10071] <= 16'hFFFF;
rommem[10072] <= 16'hFFFF;
rommem[10073] <= 16'hFFFF;
rommem[10074] <= 16'hFFFF;
rommem[10075] <= 16'hFFFF;
rommem[10076] <= 16'hFFFF;
rommem[10077] <= 16'hFFFF;
rommem[10078] <= 16'hFFFF;
rommem[10079] <= 16'hFFFF;
rommem[10080] <= 16'hFFFF;
rommem[10081] <= 16'hFFFF;
rommem[10082] <= 16'hFFFF;
rommem[10083] <= 16'hFFFF;
rommem[10084] <= 16'hFFFF;
rommem[10085] <= 16'hFFFF;
rommem[10086] <= 16'hFFFF;
rommem[10087] <= 16'hFFFF;
rommem[10088] <= 16'hFFFF;
rommem[10089] <= 16'hFFFF;
rommem[10090] <= 16'hFFFF;
rommem[10091] <= 16'hFFFF;
rommem[10092] <= 16'hFFFF;
rommem[10093] <= 16'hFFFF;
rommem[10094] <= 16'hFFFF;
rommem[10095] <= 16'hFFFF;
rommem[10096] <= 16'hFFFF;
rommem[10097] <= 16'hFFFF;
rommem[10098] <= 16'hFFFF;
rommem[10099] <= 16'hFFFF;
rommem[10100] <= 16'hFFFF;
rommem[10101] <= 16'hFFFF;
rommem[10102] <= 16'hFFFF;
rommem[10103] <= 16'hFFFF;
rommem[10104] <= 16'hFFFF;
rommem[10105] <= 16'hFFFF;
rommem[10106] <= 16'hFFFF;
rommem[10107] <= 16'hFFFF;
rommem[10108] <= 16'hFFFF;
rommem[10109] <= 16'hFFFF;
rommem[10110] <= 16'hFFFF;
rommem[10111] <= 16'hFFFF;
rommem[10112] <= 16'hFFFF;
rommem[10113] <= 16'hFFFF;
rommem[10114] <= 16'hFFFF;
rommem[10115] <= 16'hFFFF;
rommem[10116] <= 16'hFFFF;
rommem[10117] <= 16'hFFFF;
rommem[10118] <= 16'hFFFF;
rommem[10119] <= 16'hFFFF;
rommem[10120] <= 16'hFFFF;
rommem[10121] <= 16'hFFFF;
rommem[10122] <= 16'hFFFF;
rommem[10123] <= 16'hFFFF;
rommem[10124] <= 16'hFFFF;
rommem[10125] <= 16'hFFFF;
rommem[10126] <= 16'hFFFF;
rommem[10127] <= 16'hFFFF;
rommem[10128] <= 16'hFFFF;
rommem[10129] <= 16'hFFFF;
rommem[10130] <= 16'hFFFF;
rommem[10131] <= 16'hFFFF;
rommem[10132] <= 16'hFFFF;
rommem[10133] <= 16'hFFFF;
rommem[10134] <= 16'hFFFF;
rommem[10135] <= 16'hFFFF;
rommem[10136] <= 16'hFFFF;
rommem[10137] <= 16'hFFFF;
rommem[10138] <= 16'hFFFF;
rommem[10139] <= 16'hFFFF;
rommem[10140] <= 16'hFFFF;
rommem[10141] <= 16'hFFFF;
rommem[10142] <= 16'hFFFF;
rommem[10143] <= 16'hFFFF;
rommem[10144] <= 16'hFFFF;
rommem[10145] <= 16'hFFFF;
rommem[10146] <= 16'hFFFF;
rommem[10147] <= 16'hFFFF;
rommem[10148] <= 16'hFFFF;
rommem[10149] <= 16'hFFFF;
rommem[10150] <= 16'hFFFF;
rommem[10151] <= 16'hFFFF;
rommem[10152] <= 16'hFFFF;
rommem[10153] <= 16'hFFFF;
rommem[10154] <= 16'hFFFF;
rommem[10155] <= 16'hFFFF;
rommem[10156] <= 16'hFFFF;
rommem[10157] <= 16'hFFFF;
rommem[10158] <= 16'hFFFF;
rommem[10159] <= 16'hFFFF;
rommem[10160] <= 16'hFFFF;
rommem[10161] <= 16'hFFFF;
rommem[10162] <= 16'hFFFF;
rommem[10163] <= 16'hFFFF;
rommem[10164] <= 16'hFFFF;
rommem[10165] <= 16'hFFFF;
rommem[10166] <= 16'hFFFF;
rommem[10167] <= 16'hFFFF;
rommem[10168] <= 16'hFFFF;
rommem[10169] <= 16'hFFFF;
rommem[10170] <= 16'hFFFF;
rommem[10171] <= 16'hFFFF;
rommem[10172] <= 16'hFFFF;
rommem[10173] <= 16'hFFFF;
rommem[10174] <= 16'hFFFF;
rommem[10175] <= 16'hFFFF;
rommem[10176] <= 16'hFFFF;
rommem[10177] <= 16'hFFFF;
rommem[10178] <= 16'hFFFF;
rommem[10179] <= 16'hFFFF;
rommem[10180] <= 16'hFFFF;
rommem[10181] <= 16'hFFFF;
rommem[10182] <= 16'hFFFF;
rommem[10183] <= 16'hFFFF;
rommem[10184] <= 16'hFFFF;
rommem[10185] <= 16'hFFFF;
rommem[10186] <= 16'hFFFF;
rommem[10187] <= 16'hFFFF;
rommem[10188] <= 16'hFFFF;
rommem[10189] <= 16'hFFFF;
rommem[10190] <= 16'hFFFF;
rommem[10191] <= 16'hFFFF;
rommem[10192] <= 16'hFFFF;
rommem[10193] <= 16'hFFFF;
rommem[10194] <= 16'hFFFF;
rommem[10195] <= 16'hFFFF;
rommem[10196] <= 16'hFFFF;
rommem[10197] <= 16'hFFFF;
rommem[10198] <= 16'hFFFF;
rommem[10199] <= 16'hFFFF;
rommem[10200] <= 16'hFFFF;
rommem[10201] <= 16'hFFFF;
rommem[10202] <= 16'hFFFF;
rommem[10203] <= 16'hFFFF;
rommem[10204] <= 16'hFFFF;
rommem[10205] <= 16'hFFFF;
rommem[10206] <= 16'hFFFF;
rommem[10207] <= 16'hFFFF;
rommem[10208] <= 16'hFFFF;
rommem[10209] <= 16'hFFFF;
rommem[10210] <= 16'hFFFF;
rommem[10211] <= 16'hFFFF;
rommem[10212] <= 16'hFFFF;
rommem[10213] <= 16'hFFFF;
rommem[10214] <= 16'hFFFF;
rommem[10215] <= 16'hFFFF;
rommem[10216] <= 16'hFFFF;
rommem[10217] <= 16'hFFFF;
rommem[10218] <= 16'hFFFF;
rommem[10219] <= 16'hFFFF;
rommem[10220] <= 16'hFFFF;
rommem[10221] <= 16'hFFFF;
rommem[10222] <= 16'hFFFF;
rommem[10223] <= 16'hFFFF;
rommem[10224] <= 16'hFFFF;
rommem[10225] <= 16'hFFFF;
rommem[10226] <= 16'hFFFF;
rommem[10227] <= 16'hFFFF;
rommem[10228] <= 16'hFFFF;
rommem[10229] <= 16'hFFFF;
rommem[10230] <= 16'hFFFF;
rommem[10231] <= 16'hFFFF;
rommem[10232] <= 16'hFFFF;
rommem[10233] <= 16'hFFFF;
rommem[10234] <= 16'hFFFF;
rommem[10235] <= 16'hFFFF;
rommem[10236] <= 16'hFFFF;
rommem[10237] <= 16'hFFFF;
rommem[10238] <= 16'hFFFF;
rommem[10239] <= 16'hFFFF;
rommem[10240] <= 16'hFFFF;
rommem[10241] <= 16'hFFFF;
rommem[10242] <= 16'hFFFF;
rommem[10243] <= 16'hFFFF;
rommem[10244] <= 16'hFFFF;
rommem[10245] <= 16'hFFFF;
rommem[10246] <= 16'hFFFF;
rommem[10247] <= 16'hFFFF;
rommem[10248] <= 16'hFFFF;
rommem[10249] <= 16'hFFFF;
rommem[10250] <= 16'hFFFF;
rommem[10251] <= 16'hFFFF;
rommem[10252] <= 16'hFFFF;
rommem[10253] <= 16'hFFFF;
rommem[10254] <= 16'hFFFF;
rommem[10255] <= 16'hFFFF;
rommem[10256] <= 16'hFFFF;
rommem[10257] <= 16'hFFFF;
rommem[10258] <= 16'hFFFF;
rommem[10259] <= 16'hFFFF;
rommem[10260] <= 16'hFFFF;
rommem[10261] <= 16'hFFFF;
rommem[10262] <= 16'hFFFF;
rommem[10263] <= 16'hFFFF;
rommem[10264] <= 16'hFFFF;
rommem[10265] <= 16'hFFFF;
rommem[10266] <= 16'hFFFF;
rommem[10267] <= 16'hFFFF;
rommem[10268] <= 16'hFFFF;
rommem[10269] <= 16'hFFFF;
rommem[10270] <= 16'hFFFF;
rommem[10271] <= 16'hFFFF;
rommem[10272] <= 16'hFFFF;
rommem[10273] <= 16'hFFFF;
rommem[10274] <= 16'hFFFF;
rommem[10275] <= 16'hFFFF;
rommem[10276] <= 16'hFFFF;
rommem[10277] <= 16'hFFFF;
rommem[10278] <= 16'hFFFF;
rommem[10279] <= 16'hFFFF;
rommem[10280] <= 16'hFFFF;
rommem[10281] <= 16'hFFFF;
rommem[10282] <= 16'hFFFF;
rommem[10283] <= 16'hFFFF;
rommem[10284] <= 16'hFFFF;
rommem[10285] <= 16'hFFFF;
rommem[10286] <= 16'hFFFF;
rommem[10287] <= 16'hFFFF;
rommem[10288] <= 16'hFFFF;
rommem[10289] <= 16'hFFFF;
rommem[10290] <= 16'hFFFF;
rommem[10291] <= 16'hFFFF;
rommem[10292] <= 16'hFFFF;
rommem[10293] <= 16'hFFFF;
rommem[10294] <= 16'hFFFF;
rommem[10295] <= 16'hFFFF;
rommem[10296] <= 16'hFFFF;
rommem[10297] <= 16'hFFFF;
rommem[10298] <= 16'hFFFF;
rommem[10299] <= 16'hFFFF;
rommem[10300] <= 16'hFFFF;
rommem[10301] <= 16'hFFFF;
rommem[10302] <= 16'hFFFF;
rommem[10303] <= 16'hFFFF;
rommem[10304] <= 16'hFFFF;
rommem[10305] <= 16'hFFFF;
rommem[10306] <= 16'hFFFF;
rommem[10307] <= 16'hFFFF;
rommem[10308] <= 16'hFFFF;
rommem[10309] <= 16'hFFFF;
rommem[10310] <= 16'hFFFF;
rommem[10311] <= 16'hFFFF;
rommem[10312] <= 16'hFFFF;
rommem[10313] <= 16'hFFFF;
rommem[10314] <= 16'hFFFF;
rommem[10315] <= 16'hFFFF;
rommem[10316] <= 16'hFFFF;
rommem[10317] <= 16'hFFFF;
rommem[10318] <= 16'hFFFF;
rommem[10319] <= 16'hFFFF;
rommem[10320] <= 16'hFFFF;
rommem[10321] <= 16'hFFFF;
rommem[10322] <= 16'hFFFF;
rommem[10323] <= 16'hFFFF;
rommem[10324] <= 16'hFFFF;
rommem[10325] <= 16'hFFFF;
rommem[10326] <= 16'hFFFF;
rommem[10327] <= 16'hFFFF;
rommem[10328] <= 16'hFFFF;
rommem[10329] <= 16'hFFFF;
rommem[10330] <= 16'hFFFF;
rommem[10331] <= 16'hFFFF;
rommem[10332] <= 16'hFFFF;
rommem[10333] <= 16'hFFFF;
rommem[10334] <= 16'hFFFF;
rommem[10335] <= 16'hFFFF;
rommem[10336] <= 16'hFFFF;
rommem[10337] <= 16'hFFFF;
rommem[10338] <= 16'hFFFF;
rommem[10339] <= 16'hFFFF;
rommem[10340] <= 16'hFFFF;
rommem[10341] <= 16'hFFFF;
rommem[10342] <= 16'hFFFF;
rommem[10343] <= 16'hFFFF;
rommem[10344] <= 16'hFFFF;
rommem[10345] <= 16'hFFFF;
rommem[10346] <= 16'hFFFF;
rommem[10347] <= 16'hFFFF;
rommem[10348] <= 16'hFFFF;
rommem[10349] <= 16'hFFFF;
rommem[10350] <= 16'hFFFF;
rommem[10351] <= 16'hFFFF;
rommem[10352] <= 16'hFFFF;
rommem[10353] <= 16'hFFFF;
rommem[10354] <= 16'hFFFF;
rommem[10355] <= 16'hFFFF;
rommem[10356] <= 16'hFFFF;
rommem[10357] <= 16'hFFFF;
rommem[10358] <= 16'hFFFF;
rommem[10359] <= 16'hFFFF;
rommem[10360] <= 16'hFFFF;
rommem[10361] <= 16'hFFFF;
rommem[10362] <= 16'hFFFF;
rommem[10363] <= 16'hFFFF;
rommem[10364] <= 16'hFFFF;
rommem[10365] <= 16'hFFFF;
rommem[10366] <= 16'hFFFF;
rommem[10367] <= 16'hFFFF;
rommem[10368] <= 16'hFFFF;
rommem[10369] <= 16'hFFFF;
rommem[10370] <= 16'hFFFF;
rommem[10371] <= 16'hFFFF;
rommem[10372] <= 16'hFFFF;
rommem[10373] <= 16'hFFFF;
rommem[10374] <= 16'hFFFF;
rommem[10375] <= 16'hFFFF;
rommem[10376] <= 16'hFFFF;
rommem[10377] <= 16'hFFFF;
rommem[10378] <= 16'hFFFF;
rommem[10379] <= 16'hFFFF;
rommem[10380] <= 16'hFFFF;
rommem[10381] <= 16'hFFFF;
rommem[10382] <= 16'hFFFF;
rommem[10383] <= 16'hFFFF;
rommem[10384] <= 16'hFFFF;
rommem[10385] <= 16'hFFFF;
rommem[10386] <= 16'hFFFF;
rommem[10387] <= 16'hFFFF;
rommem[10388] <= 16'hFFFF;
rommem[10389] <= 16'hFFFF;
rommem[10390] <= 16'hFFFF;
rommem[10391] <= 16'hFFFF;
rommem[10392] <= 16'hFFFF;
rommem[10393] <= 16'hFFFF;
rommem[10394] <= 16'hFFFF;
rommem[10395] <= 16'hFFFF;
rommem[10396] <= 16'hFFFF;
rommem[10397] <= 16'hFFFF;
rommem[10398] <= 16'hFFFF;
rommem[10399] <= 16'hFFFF;
rommem[10400] <= 16'hFFFF;
rommem[10401] <= 16'hFFFF;
rommem[10402] <= 16'hFFFF;
rommem[10403] <= 16'hFFFF;
rommem[10404] <= 16'hFFFF;
rommem[10405] <= 16'hFFFF;
rommem[10406] <= 16'hFFFF;
rommem[10407] <= 16'hFFFF;
rommem[10408] <= 16'hFFFF;
rommem[10409] <= 16'hFFFF;
rommem[10410] <= 16'hFFFF;
rommem[10411] <= 16'hFFFF;
rommem[10412] <= 16'hFFFF;
rommem[10413] <= 16'hFFFF;
rommem[10414] <= 16'hFFFF;
rommem[10415] <= 16'hFFFF;
rommem[10416] <= 16'hFFFF;
rommem[10417] <= 16'hFFFF;
rommem[10418] <= 16'hFFFF;
rommem[10419] <= 16'hFFFF;
rommem[10420] <= 16'hFFFF;
rommem[10421] <= 16'hFFFF;
rommem[10422] <= 16'hFFFF;
rommem[10423] <= 16'hFFFF;
rommem[10424] <= 16'hFFFF;
rommem[10425] <= 16'hFFFF;
rommem[10426] <= 16'hFFFF;
rommem[10427] <= 16'hFFFF;
rommem[10428] <= 16'hFFFF;
rommem[10429] <= 16'hFFFF;
rommem[10430] <= 16'hFFFF;
rommem[10431] <= 16'hFFFF;
rommem[10432] <= 16'hFFFF;
rommem[10433] <= 16'hFFFF;
rommem[10434] <= 16'hFFFF;
rommem[10435] <= 16'hFFFF;
rommem[10436] <= 16'hFFFF;
rommem[10437] <= 16'hFFFF;
rommem[10438] <= 16'hFFFF;
rommem[10439] <= 16'hFFFF;
rommem[10440] <= 16'hFFFF;
rommem[10441] <= 16'hFFFF;
rommem[10442] <= 16'hFFFF;
rommem[10443] <= 16'hFFFF;
rommem[10444] <= 16'hFFFF;
rommem[10445] <= 16'hFFFF;
rommem[10446] <= 16'hFFFF;
rommem[10447] <= 16'hFFFF;
rommem[10448] <= 16'hFFFF;
rommem[10449] <= 16'hFFFF;
rommem[10450] <= 16'hFFFF;
rommem[10451] <= 16'hFFFF;
rommem[10452] <= 16'hFFFF;
rommem[10453] <= 16'hFFFF;
rommem[10454] <= 16'hFFFF;
rommem[10455] <= 16'hFFFF;
rommem[10456] <= 16'hFFFF;
rommem[10457] <= 16'hFFFF;
rommem[10458] <= 16'hFFFF;
rommem[10459] <= 16'hFFFF;
rommem[10460] <= 16'hFFFF;
rommem[10461] <= 16'hFFFF;
rommem[10462] <= 16'hFFFF;
rommem[10463] <= 16'hFFFF;
rommem[10464] <= 16'hFFFF;
rommem[10465] <= 16'hFFFF;
rommem[10466] <= 16'hFFFF;
rommem[10467] <= 16'hFFFF;
rommem[10468] <= 16'hFFFF;
rommem[10469] <= 16'hFFFF;
rommem[10470] <= 16'hFFFF;
rommem[10471] <= 16'hFFFF;
rommem[10472] <= 16'hFFFF;
rommem[10473] <= 16'hFFFF;
rommem[10474] <= 16'hFFFF;
rommem[10475] <= 16'hFFFF;
rommem[10476] <= 16'hFFFF;
rommem[10477] <= 16'hFFFF;
rommem[10478] <= 16'hFFFF;
rommem[10479] <= 16'hFFFF;
rommem[10480] <= 16'hFFFF;
rommem[10481] <= 16'hFFFF;
rommem[10482] <= 16'hFFFF;
rommem[10483] <= 16'hFFFF;
rommem[10484] <= 16'hFFFF;
rommem[10485] <= 16'hFFFF;
rommem[10486] <= 16'hFFFF;
rommem[10487] <= 16'hFFFF;
rommem[10488] <= 16'hFFFF;
rommem[10489] <= 16'hFFFF;
rommem[10490] <= 16'hFFFF;
rommem[10491] <= 16'hFFFF;
rommem[10492] <= 16'hFFFF;
rommem[10493] <= 16'hFFFF;
rommem[10494] <= 16'hFFFF;
rommem[10495] <= 16'hFFFF;
rommem[10496] <= 16'hFFFF;
rommem[10497] <= 16'hFFFF;
rommem[10498] <= 16'hFFFF;
rommem[10499] <= 16'hFFFF;
rommem[10500] <= 16'hFFFF;
rommem[10501] <= 16'hFFFF;
rommem[10502] <= 16'hFFFF;
rommem[10503] <= 16'hFFFF;
rommem[10504] <= 16'hFFFF;
rommem[10505] <= 16'hFFFF;
rommem[10506] <= 16'hFFFF;
rommem[10507] <= 16'hFFFF;
rommem[10508] <= 16'hFFFF;
rommem[10509] <= 16'hFFFF;
rommem[10510] <= 16'hFFFF;
rommem[10511] <= 16'hFFFF;
rommem[10512] <= 16'hFFFF;
rommem[10513] <= 16'hFFFF;
rommem[10514] <= 16'hFFFF;
rommem[10515] <= 16'hFFFF;
rommem[10516] <= 16'hFFFF;
rommem[10517] <= 16'hFFFF;
rommem[10518] <= 16'hFFFF;
rommem[10519] <= 16'hFFFF;
rommem[10520] <= 16'hFFFF;
rommem[10521] <= 16'hFFFF;
rommem[10522] <= 16'hFFFF;
rommem[10523] <= 16'hFFFF;
rommem[10524] <= 16'hFFFF;
rommem[10525] <= 16'hFFFF;
rommem[10526] <= 16'hFFFF;
rommem[10527] <= 16'hFFFF;
rommem[10528] <= 16'hFFFF;
rommem[10529] <= 16'hFFFF;
rommem[10530] <= 16'hFFFF;
rommem[10531] <= 16'hFFFF;
rommem[10532] <= 16'hFFFF;
rommem[10533] <= 16'hFFFF;
rommem[10534] <= 16'hFFFF;
rommem[10535] <= 16'hFFFF;
rommem[10536] <= 16'hFFFF;
rommem[10537] <= 16'hFFFF;
rommem[10538] <= 16'hFFFF;
rommem[10539] <= 16'hFFFF;
rommem[10540] <= 16'hFFFF;
rommem[10541] <= 16'hFFFF;
rommem[10542] <= 16'hFFFF;
rommem[10543] <= 16'hFFFF;
rommem[10544] <= 16'hFFFF;
rommem[10545] <= 16'hFFFF;
rommem[10546] <= 16'hFFFF;
rommem[10547] <= 16'hFFFF;
rommem[10548] <= 16'hFFFF;
rommem[10549] <= 16'hFFFF;
rommem[10550] <= 16'hFFFF;
rommem[10551] <= 16'hFFFF;
rommem[10552] <= 16'hFFFF;
rommem[10553] <= 16'hFFFF;
rommem[10554] <= 16'hFFFF;
rommem[10555] <= 16'hFFFF;
rommem[10556] <= 16'hFFFF;
rommem[10557] <= 16'hFFFF;
rommem[10558] <= 16'hFFFF;
rommem[10559] <= 16'hFFFF;
rommem[10560] <= 16'hFFFF;
rommem[10561] <= 16'hFFFF;
rommem[10562] <= 16'hFFFF;
rommem[10563] <= 16'hFFFF;
rommem[10564] <= 16'hFFFF;
rommem[10565] <= 16'hFFFF;
rommem[10566] <= 16'hFFFF;
rommem[10567] <= 16'hFFFF;
rommem[10568] <= 16'hFFFF;
rommem[10569] <= 16'hFFFF;
rommem[10570] <= 16'hFFFF;
rommem[10571] <= 16'hFFFF;
rommem[10572] <= 16'hFFFF;
rommem[10573] <= 16'hFFFF;
rommem[10574] <= 16'hFFFF;
rommem[10575] <= 16'hFFFF;
rommem[10576] <= 16'hFFFF;
rommem[10577] <= 16'hFFFF;
rommem[10578] <= 16'hFFFF;
rommem[10579] <= 16'hFFFF;
rommem[10580] <= 16'hFFFF;
rommem[10581] <= 16'hFFFF;
rommem[10582] <= 16'hFFFF;
rommem[10583] <= 16'hFFFF;
rommem[10584] <= 16'hFFFF;
rommem[10585] <= 16'hFFFF;
rommem[10586] <= 16'hFFFF;
rommem[10587] <= 16'hFFFF;
rommem[10588] <= 16'hFFFF;
rommem[10589] <= 16'hFFFF;
rommem[10590] <= 16'hFFFF;
rommem[10591] <= 16'hFFFF;
rommem[10592] <= 16'hFFFF;
rommem[10593] <= 16'hFFFF;
rommem[10594] <= 16'hFFFF;
rommem[10595] <= 16'hFFFF;
rommem[10596] <= 16'hFFFF;
rommem[10597] <= 16'hFFFF;
rommem[10598] <= 16'hFFFF;
rommem[10599] <= 16'hFFFF;
rommem[10600] <= 16'hFFFF;
rommem[10601] <= 16'hFFFF;
rommem[10602] <= 16'hFFFF;
rommem[10603] <= 16'hFFFF;
rommem[10604] <= 16'hFFFF;
rommem[10605] <= 16'hFFFF;
rommem[10606] <= 16'hFFFF;
rommem[10607] <= 16'hFFFF;
rommem[10608] <= 16'hFFFF;
rommem[10609] <= 16'hFFFF;
rommem[10610] <= 16'hFFFF;
rommem[10611] <= 16'hFFFF;
rommem[10612] <= 16'hFFFF;
rommem[10613] <= 16'hFFFF;
rommem[10614] <= 16'hFFFF;
rommem[10615] <= 16'hFFFF;
rommem[10616] <= 16'hFFFF;
rommem[10617] <= 16'hFFFF;
rommem[10618] <= 16'hFFFF;
rommem[10619] <= 16'hFFFF;
rommem[10620] <= 16'hFFFF;
rommem[10621] <= 16'hFFFF;
rommem[10622] <= 16'hFFFF;
rommem[10623] <= 16'hFFFF;
rommem[10624] <= 16'hFFFF;
rommem[10625] <= 16'hFFFF;
rommem[10626] <= 16'hFFFF;
rommem[10627] <= 16'hFFFF;
rommem[10628] <= 16'hFFFF;
rommem[10629] <= 16'hFFFF;
rommem[10630] <= 16'hFFFF;
rommem[10631] <= 16'hFFFF;
rommem[10632] <= 16'hFFFF;
rommem[10633] <= 16'hFFFF;
rommem[10634] <= 16'hFFFF;
rommem[10635] <= 16'hFFFF;
rommem[10636] <= 16'hFFFF;
rommem[10637] <= 16'hFFFF;
rommem[10638] <= 16'hFFFF;
rommem[10639] <= 16'hFFFF;
rommem[10640] <= 16'hFFFF;
rommem[10641] <= 16'hFFFF;
rommem[10642] <= 16'hFFFF;
rommem[10643] <= 16'hFFFF;
rommem[10644] <= 16'hFFFF;
rommem[10645] <= 16'hFFFF;
rommem[10646] <= 16'hFFFF;
rommem[10647] <= 16'hFFFF;
rommem[10648] <= 16'hFFFF;
rommem[10649] <= 16'hFFFF;
rommem[10650] <= 16'hFFFF;
rommem[10651] <= 16'hFFFF;
rommem[10652] <= 16'hFFFF;
rommem[10653] <= 16'hFFFF;
rommem[10654] <= 16'hFFFF;
rommem[10655] <= 16'hFFFF;
rommem[10656] <= 16'hFFFF;
rommem[10657] <= 16'hFFFF;
rommem[10658] <= 16'hFFFF;
rommem[10659] <= 16'hFFFF;
rommem[10660] <= 16'hFFFF;
rommem[10661] <= 16'hFFFF;
rommem[10662] <= 16'hFFFF;
rommem[10663] <= 16'hFFFF;
rommem[10664] <= 16'hFFFF;
rommem[10665] <= 16'hFFFF;
rommem[10666] <= 16'hFFFF;
rommem[10667] <= 16'hFFFF;
rommem[10668] <= 16'hFFFF;
rommem[10669] <= 16'hFFFF;
rommem[10670] <= 16'hFFFF;
rommem[10671] <= 16'hFFFF;
rommem[10672] <= 16'hFFFF;
rommem[10673] <= 16'hFFFF;
rommem[10674] <= 16'hFFFF;
rommem[10675] <= 16'hFFFF;
rommem[10676] <= 16'hFFFF;
rommem[10677] <= 16'hFFFF;
rommem[10678] <= 16'hFFFF;
rommem[10679] <= 16'hFFFF;
rommem[10680] <= 16'hFFFF;
rommem[10681] <= 16'hFFFF;
rommem[10682] <= 16'hFFFF;
rommem[10683] <= 16'hFFFF;
rommem[10684] <= 16'hFFFF;
rommem[10685] <= 16'hFFFF;
rommem[10686] <= 16'hFFFF;
rommem[10687] <= 16'hFFFF;
rommem[10688] <= 16'hFFFF;
rommem[10689] <= 16'hFFFF;
rommem[10690] <= 16'hFFFF;
rommem[10691] <= 16'hFFFF;
rommem[10692] <= 16'hFFFF;
rommem[10693] <= 16'hFFFF;
rommem[10694] <= 16'hFFFF;
rommem[10695] <= 16'hFFFF;
rommem[10696] <= 16'hFFFF;
rommem[10697] <= 16'hFFFF;
rommem[10698] <= 16'hFFFF;
rommem[10699] <= 16'hFFFF;
rommem[10700] <= 16'hFFFF;
rommem[10701] <= 16'hFFFF;
rommem[10702] <= 16'hFFFF;
rommem[10703] <= 16'hFFFF;
rommem[10704] <= 16'hFFFF;
rommem[10705] <= 16'hFFFF;
rommem[10706] <= 16'hFFFF;
rommem[10707] <= 16'hFFFF;
rommem[10708] <= 16'hFFFF;
rommem[10709] <= 16'hFFFF;
rommem[10710] <= 16'hFFFF;
rommem[10711] <= 16'hFFFF;
rommem[10712] <= 16'hFFFF;
rommem[10713] <= 16'hFFFF;
rommem[10714] <= 16'hFFFF;
rommem[10715] <= 16'hFFFF;
rommem[10716] <= 16'hFFFF;
rommem[10717] <= 16'hFFFF;
rommem[10718] <= 16'hFFFF;
rommem[10719] <= 16'hFFFF;
rommem[10720] <= 16'hFFFF;
rommem[10721] <= 16'hFFFF;
rommem[10722] <= 16'hFFFF;
rommem[10723] <= 16'hFFFF;
rommem[10724] <= 16'hFFFF;
rommem[10725] <= 16'hFFFF;
rommem[10726] <= 16'hFFFF;
rommem[10727] <= 16'hFFFF;
rommem[10728] <= 16'hFFFF;
rommem[10729] <= 16'hFFFF;
rommem[10730] <= 16'hFFFF;
rommem[10731] <= 16'hFFFF;
rommem[10732] <= 16'hFFFF;
rommem[10733] <= 16'hFFFF;
rommem[10734] <= 16'hFFFF;
rommem[10735] <= 16'hFFFF;
rommem[10736] <= 16'hFFFF;
rommem[10737] <= 16'hFFFF;
rommem[10738] <= 16'hFFFF;
rommem[10739] <= 16'hFFFF;
rommem[10740] <= 16'hFFFF;
rommem[10741] <= 16'hFFFF;
rommem[10742] <= 16'hFFFF;
rommem[10743] <= 16'hFFFF;
rommem[10744] <= 16'hFFFF;
rommem[10745] <= 16'hFFFF;
rommem[10746] <= 16'hFFFF;
rommem[10747] <= 16'hFFFF;
rommem[10748] <= 16'hFFFF;
rommem[10749] <= 16'hFFFF;
rommem[10750] <= 16'hFFFF;
rommem[10751] <= 16'hFFFF;
rommem[10752] <= 16'hFFFF;
rommem[10753] <= 16'hFFFF;
rommem[10754] <= 16'hFFFF;
rommem[10755] <= 16'hFFFF;
rommem[10756] <= 16'hFFFF;
rommem[10757] <= 16'hFFFF;
rommem[10758] <= 16'hFFFF;
rommem[10759] <= 16'hFFFF;
rommem[10760] <= 16'hFFFF;
rommem[10761] <= 16'hFFFF;
rommem[10762] <= 16'hFFFF;
rommem[10763] <= 16'hFFFF;
rommem[10764] <= 16'hFFFF;
rommem[10765] <= 16'hFFFF;
rommem[10766] <= 16'hFFFF;
rommem[10767] <= 16'hFFFF;
rommem[10768] <= 16'hFFFF;
rommem[10769] <= 16'hFFFF;
rommem[10770] <= 16'hFFFF;
rommem[10771] <= 16'hFFFF;
rommem[10772] <= 16'hFFFF;
rommem[10773] <= 16'hFFFF;
rommem[10774] <= 16'hFFFF;
rommem[10775] <= 16'hFFFF;
rommem[10776] <= 16'hFFFF;
rommem[10777] <= 16'hFFFF;
rommem[10778] <= 16'hFFFF;
rommem[10779] <= 16'hFFFF;
rommem[10780] <= 16'hFFFF;
rommem[10781] <= 16'hFFFF;
rommem[10782] <= 16'hFFFF;
rommem[10783] <= 16'hFFFF;
rommem[10784] <= 16'hFFFF;
rommem[10785] <= 16'hFFFF;
rommem[10786] <= 16'hFFFF;
rommem[10787] <= 16'hFFFF;
rommem[10788] <= 16'hFFFF;
rommem[10789] <= 16'hFFFF;
rommem[10790] <= 16'hFFFF;
rommem[10791] <= 16'hFFFF;
rommem[10792] <= 16'hFFFF;
rommem[10793] <= 16'hFFFF;
rommem[10794] <= 16'hFFFF;
rommem[10795] <= 16'hFFFF;
rommem[10796] <= 16'hFFFF;
rommem[10797] <= 16'hFFFF;
rommem[10798] <= 16'hFFFF;
rommem[10799] <= 16'hFFFF;
rommem[10800] <= 16'hFFFF;
rommem[10801] <= 16'hFFFF;
rommem[10802] <= 16'hFFFF;
rommem[10803] <= 16'hFFFF;
rommem[10804] <= 16'hFFFF;
rommem[10805] <= 16'hFFFF;
rommem[10806] <= 16'hFFFF;
rommem[10807] <= 16'hFFFF;
rommem[10808] <= 16'hFFFF;
rommem[10809] <= 16'hFFFF;
rommem[10810] <= 16'hFFFF;
rommem[10811] <= 16'hFFFF;
rommem[10812] <= 16'hFFFF;
rommem[10813] <= 16'hFFFF;
rommem[10814] <= 16'hFFFF;
rommem[10815] <= 16'hFFFF;
rommem[10816] <= 16'hFFFF;
rommem[10817] <= 16'hFFFF;
rommem[10818] <= 16'hFFFF;
rommem[10819] <= 16'hFFFF;
rommem[10820] <= 16'hFFFF;
rommem[10821] <= 16'hFFFF;
rommem[10822] <= 16'hFFFF;
rommem[10823] <= 16'hFFFF;
rommem[10824] <= 16'hFFFF;
rommem[10825] <= 16'hFFFF;
rommem[10826] <= 16'hFFFF;
rommem[10827] <= 16'hFFFF;
rommem[10828] <= 16'hFFFF;
rommem[10829] <= 16'hFFFF;
rommem[10830] <= 16'hFFFF;
rommem[10831] <= 16'hFFFF;
rommem[10832] <= 16'hFFFF;
rommem[10833] <= 16'hFFFF;
rommem[10834] <= 16'hFFFF;
rommem[10835] <= 16'hFFFF;
rommem[10836] <= 16'hFFFF;
rommem[10837] <= 16'hFFFF;
rommem[10838] <= 16'hFFFF;
rommem[10839] <= 16'hFFFF;
rommem[10840] <= 16'hFFFF;
rommem[10841] <= 16'hFFFF;
rommem[10842] <= 16'hFFFF;
rommem[10843] <= 16'hFFFF;
rommem[10844] <= 16'hFFFF;
rommem[10845] <= 16'hFFFF;
rommem[10846] <= 16'hFFFF;
rommem[10847] <= 16'hFFFF;
rommem[10848] <= 16'hFFFF;
rommem[10849] <= 16'hFFFF;
rommem[10850] <= 16'hFFFF;
rommem[10851] <= 16'hFFFF;
rommem[10852] <= 16'hFFFF;
rommem[10853] <= 16'hFFFF;
rommem[10854] <= 16'hFFFF;
rommem[10855] <= 16'hFFFF;
rommem[10856] <= 16'hFFFF;
rommem[10857] <= 16'hFFFF;
rommem[10858] <= 16'hFFFF;
rommem[10859] <= 16'hFFFF;
rommem[10860] <= 16'hFFFF;
rommem[10861] <= 16'hFFFF;
rommem[10862] <= 16'hFFFF;
rommem[10863] <= 16'hFFFF;
rommem[10864] <= 16'hFFFF;
rommem[10865] <= 16'hFFFF;
rommem[10866] <= 16'hFFFF;
rommem[10867] <= 16'hFFFF;
rommem[10868] <= 16'hFFFF;
rommem[10869] <= 16'hFFFF;
rommem[10870] <= 16'hFFFF;
rommem[10871] <= 16'hFFFF;
rommem[10872] <= 16'hFFFF;
rommem[10873] <= 16'hFFFF;
rommem[10874] <= 16'hFFFF;
rommem[10875] <= 16'hFFFF;
rommem[10876] <= 16'hFFFF;
rommem[10877] <= 16'hFFFF;
rommem[10878] <= 16'hFFFF;
rommem[10879] <= 16'hFFFF;
rommem[10880] <= 16'hFFFF;
rommem[10881] <= 16'hFFFF;
rommem[10882] <= 16'hFFFF;
rommem[10883] <= 16'hFFFF;
rommem[10884] <= 16'hFFFF;
rommem[10885] <= 16'hFFFF;
rommem[10886] <= 16'hFFFF;
rommem[10887] <= 16'hFFFF;
rommem[10888] <= 16'hFFFF;
rommem[10889] <= 16'hFFFF;
rommem[10890] <= 16'hFFFF;
rommem[10891] <= 16'hFFFF;
rommem[10892] <= 16'hFFFF;
rommem[10893] <= 16'hFFFF;
rommem[10894] <= 16'hFFFF;
rommem[10895] <= 16'hFFFF;
rommem[10896] <= 16'hFFFF;
rommem[10897] <= 16'hFFFF;
rommem[10898] <= 16'hFFFF;
rommem[10899] <= 16'hFFFF;
rommem[10900] <= 16'hFFFF;
rommem[10901] <= 16'hFFFF;
rommem[10902] <= 16'hFFFF;
rommem[10903] <= 16'hFFFF;
rommem[10904] <= 16'hFFFF;
rommem[10905] <= 16'hFFFF;
rommem[10906] <= 16'hFFFF;
rommem[10907] <= 16'hFFFF;
rommem[10908] <= 16'hFFFF;
rommem[10909] <= 16'hFFFF;
rommem[10910] <= 16'hFFFF;
rommem[10911] <= 16'hFFFF;
rommem[10912] <= 16'hFFFF;
rommem[10913] <= 16'hFFFF;
rommem[10914] <= 16'hFFFF;
rommem[10915] <= 16'hFFFF;
rommem[10916] <= 16'hFFFF;
rommem[10917] <= 16'hFFFF;
rommem[10918] <= 16'hFFFF;
rommem[10919] <= 16'hFFFF;
rommem[10920] <= 16'hFFFF;
rommem[10921] <= 16'hFFFF;
rommem[10922] <= 16'hFFFF;
rommem[10923] <= 16'hFFFF;
rommem[10924] <= 16'hFFFF;
rommem[10925] <= 16'hFFFF;
rommem[10926] <= 16'hFFFF;
rommem[10927] <= 16'hFFFF;
rommem[10928] <= 16'hFFFF;
rommem[10929] <= 16'hFFFF;
rommem[10930] <= 16'hFFFF;
rommem[10931] <= 16'hFFFF;
rommem[10932] <= 16'hFFFF;
rommem[10933] <= 16'hFFFF;
rommem[10934] <= 16'hFFFF;
rommem[10935] <= 16'hFFFF;
rommem[10936] <= 16'hFFFF;
rommem[10937] <= 16'hFFFF;
rommem[10938] <= 16'hFFFF;
rommem[10939] <= 16'hFFFF;
rommem[10940] <= 16'hFFFF;
rommem[10941] <= 16'hFFFF;
rommem[10942] <= 16'hFFFF;
rommem[10943] <= 16'hFFFF;
rommem[10944] <= 16'hFFFF;
rommem[10945] <= 16'hFFFF;
rommem[10946] <= 16'hFFFF;
rommem[10947] <= 16'hFFFF;
rommem[10948] <= 16'hFFFF;
rommem[10949] <= 16'hFFFF;
rommem[10950] <= 16'hFFFF;
rommem[10951] <= 16'hFFFF;
rommem[10952] <= 16'hFFFF;
rommem[10953] <= 16'hFFFF;
rommem[10954] <= 16'hFFFF;
rommem[10955] <= 16'hFFFF;
rommem[10956] <= 16'hFFFF;
rommem[10957] <= 16'hFFFF;
rommem[10958] <= 16'hFFFF;
rommem[10959] <= 16'hFFFF;
rommem[10960] <= 16'hFFFF;
rommem[10961] <= 16'hFFFF;
rommem[10962] <= 16'hFFFF;
rommem[10963] <= 16'hFFFF;
rommem[10964] <= 16'hFFFF;
rommem[10965] <= 16'hFFFF;
rommem[10966] <= 16'hFFFF;
rommem[10967] <= 16'hFFFF;
rommem[10968] <= 16'hFFFF;
rommem[10969] <= 16'hFFFF;
rommem[10970] <= 16'hFFFF;
rommem[10971] <= 16'hFFFF;
rommem[10972] <= 16'hFFFF;
rommem[10973] <= 16'hFFFF;
rommem[10974] <= 16'hFFFF;
rommem[10975] <= 16'hFFFF;
rommem[10976] <= 16'hFFFF;
rommem[10977] <= 16'hFFFF;
rommem[10978] <= 16'hFFFF;
rommem[10979] <= 16'hFFFF;
rommem[10980] <= 16'hFFFF;
rommem[10981] <= 16'hFFFF;
rommem[10982] <= 16'hFFFF;
rommem[10983] <= 16'hFFFF;
rommem[10984] <= 16'hFFFF;
rommem[10985] <= 16'hFFFF;
rommem[10986] <= 16'hFFFF;
rommem[10987] <= 16'hFFFF;
rommem[10988] <= 16'hFFFF;
rommem[10989] <= 16'hFFFF;
rommem[10990] <= 16'hFFFF;
rommem[10991] <= 16'hFFFF;
rommem[10992] <= 16'hFFFF;
rommem[10993] <= 16'hFFFF;
rommem[10994] <= 16'hFFFF;
rommem[10995] <= 16'hFFFF;
rommem[10996] <= 16'hFFFF;
rommem[10997] <= 16'hFFFF;
rommem[10998] <= 16'hFFFF;
rommem[10999] <= 16'hFFFF;
rommem[11000] <= 16'hFFFF;
rommem[11001] <= 16'hFFFF;
rommem[11002] <= 16'hFFFF;
rommem[11003] <= 16'hFFFF;
rommem[11004] <= 16'hFFFF;
rommem[11005] <= 16'hFFFF;
rommem[11006] <= 16'hFFFF;
rommem[11007] <= 16'hFFFF;
rommem[11008] <= 16'hFFFF;
rommem[11009] <= 16'hFFFF;
rommem[11010] <= 16'hFFFF;
rommem[11011] <= 16'hFFFF;
rommem[11012] <= 16'hFFFF;
rommem[11013] <= 16'hFFFF;
rommem[11014] <= 16'hFFFF;
rommem[11015] <= 16'hFFFF;
rommem[11016] <= 16'hFFFF;
rommem[11017] <= 16'hFFFF;
rommem[11018] <= 16'hFFFF;
rommem[11019] <= 16'hFFFF;
rommem[11020] <= 16'hFFFF;
rommem[11021] <= 16'hFFFF;
rommem[11022] <= 16'hFFFF;
rommem[11023] <= 16'hFFFF;
rommem[11024] <= 16'hFFFF;
rommem[11025] <= 16'hFFFF;
rommem[11026] <= 16'hFFFF;
rommem[11027] <= 16'hFFFF;
rommem[11028] <= 16'hFFFF;
rommem[11029] <= 16'hFFFF;
rommem[11030] <= 16'hFFFF;
rommem[11031] <= 16'hFFFF;
rommem[11032] <= 16'hFFFF;
rommem[11033] <= 16'hFFFF;
rommem[11034] <= 16'hFFFF;
rommem[11035] <= 16'hFFFF;
rommem[11036] <= 16'hFFFF;
rommem[11037] <= 16'hFFFF;
rommem[11038] <= 16'hFFFF;
rommem[11039] <= 16'hFFFF;
rommem[11040] <= 16'hFFFF;
rommem[11041] <= 16'hFFFF;
rommem[11042] <= 16'hFFFF;
rommem[11043] <= 16'hFFFF;
rommem[11044] <= 16'hFFFF;
rommem[11045] <= 16'hFFFF;
rommem[11046] <= 16'hFFFF;
rommem[11047] <= 16'hFFFF;
rommem[11048] <= 16'hFFFF;
rommem[11049] <= 16'hFFFF;
rommem[11050] <= 16'hFFFF;
rommem[11051] <= 16'hFFFF;
rommem[11052] <= 16'hFFFF;
rommem[11053] <= 16'hFFFF;
rommem[11054] <= 16'hFFFF;
rommem[11055] <= 16'hFFFF;
rommem[11056] <= 16'hFFFF;
rommem[11057] <= 16'hFFFF;
rommem[11058] <= 16'hFFFF;
rommem[11059] <= 16'hFFFF;
rommem[11060] <= 16'hFFFF;
rommem[11061] <= 16'hFFFF;
rommem[11062] <= 16'hFFFF;
rommem[11063] <= 16'hFFFF;
rommem[11064] <= 16'hFFFF;
rommem[11065] <= 16'hFFFF;
rommem[11066] <= 16'hFFFF;
rommem[11067] <= 16'hFFFF;
rommem[11068] <= 16'hFFFF;
rommem[11069] <= 16'hFFFF;
rommem[11070] <= 16'hFFFF;
rommem[11071] <= 16'hFFFF;
rommem[11072] <= 16'hFFFF;
rommem[11073] <= 16'hFFFF;
rommem[11074] <= 16'hFFFF;
rommem[11075] <= 16'hFFFF;
rommem[11076] <= 16'hFFFF;
rommem[11077] <= 16'hFFFF;
rommem[11078] <= 16'hFFFF;
rommem[11079] <= 16'hFFFF;
rommem[11080] <= 16'hFFFF;
rommem[11081] <= 16'hFFFF;
rommem[11082] <= 16'hFFFF;
rommem[11083] <= 16'hFFFF;
rommem[11084] <= 16'hFFFF;
rommem[11085] <= 16'hFFFF;
rommem[11086] <= 16'hFFFF;
rommem[11087] <= 16'hFFFF;
rommem[11088] <= 16'hFFFF;
rommem[11089] <= 16'hFFFF;
rommem[11090] <= 16'hFFFF;
rommem[11091] <= 16'hFFFF;
rommem[11092] <= 16'hFFFF;
rommem[11093] <= 16'hFFFF;
rommem[11094] <= 16'hFFFF;
rommem[11095] <= 16'hFFFF;
rommem[11096] <= 16'hFFFF;
rommem[11097] <= 16'hFFFF;
rommem[11098] <= 16'hFFFF;
rommem[11099] <= 16'hFFFF;
rommem[11100] <= 16'hFFFF;
rommem[11101] <= 16'hFFFF;
rommem[11102] <= 16'hFFFF;
rommem[11103] <= 16'hFFFF;
rommem[11104] <= 16'hFFFF;
rommem[11105] <= 16'hFFFF;
rommem[11106] <= 16'hFFFF;
rommem[11107] <= 16'hFFFF;
rommem[11108] <= 16'hFFFF;
rommem[11109] <= 16'hFFFF;
rommem[11110] <= 16'hFFFF;
rommem[11111] <= 16'hFFFF;
rommem[11112] <= 16'hFFFF;
rommem[11113] <= 16'hFFFF;
rommem[11114] <= 16'hFFFF;
rommem[11115] <= 16'hFFFF;
rommem[11116] <= 16'hFFFF;
rommem[11117] <= 16'hFFFF;
rommem[11118] <= 16'hFFFF;
rommem[11119] <= 16'hFFFF;
rommem[11120] <= 16'hFFFF;
rommem[11121] <= 16'hFFFF;
rommem[11122] <= 16'hFFFF;
rommem[11123] <= 16'hFFFF;
rommem[11124] <= 16'hFFFF;
rommem[11125] <= 16'hFFFF;
rommem[11126] <= 16'hFFFF;
rommem[11127] <= 16'hFFFF;
rommem[11128] <= 16'hFFFF;
rommem[11129] <= 16'hFFFF;
rommem[11130] <= 16'hFFFF;
rommem[11131] <= 16'hFFFF;
rommem[11132] <= 16'hFFFF;
rommem[11133] <= 16'hFFFF;
rommem[11134] <= 16'hFFFF;
rommem[11135] <= 16'hFFFF;
rommem[11136] <= 16'hFFFF;
rommem[11137] <= 16'hFFFF;
rommem[11138] <= 16'hFFFF;
rommem[11139] <= 16'hFFFF;
rommem[11140] <= 16'hFFFF;
rommem[11141] <= 16'hFFFF;
rommem[11142] <= 16'hFFFF;
rommem[11143] <= 16'hFFFF;
rommem[11144] <= 16'hFFFF;
rommem[11145] <= 16'hFFFF;
rommem[11146] <= 16'hFFFF;
rommem[11147] <= 16'hFFFF;
rommem[11148] <= 16'hFFFF;
rommem[11149] <= 16'hFFFF;
rommem[11150] <= 16'hFFFF;
rommem[11151] <= 16'hFFFF;
rommem[11152] <= 16'hFFFF;
rommem[11153] <= 16'hFFFF;
rommem[11154] <= 16'hFFFF;
rommem[11155] <= 16'hFFFF;
rommem[11156] <= 16'hFFFF;
rommem[11157] <= 16'hFFFF;
rommem[11158] <= 16'hFFFF;
rommem[11159] <= 16'hFFFF;
rommem[11160] <= 16'hFFFF;
rommem[11161] <= 16'hFFFF;
rommem[11162] <= 16'hFFFF;
rommem[11163] <= 16'hFFFF;
rommem[11164] <= 16'hFFFF;
rommem[11165] <= 16'hFFFF;
rommem[11166] <= 16'hFFFF;
rommem[11167] <= 16'hFFFF;
rommem[11168] <= 16'hFFFF;
rommem[11169] <= 16'hFFFF;
rommem[11170] <= 16'hFFFF;
rommem[11171] <= 16'hFFFF;
rommem[11172] <= 16'hFFFF;
rommem[11173] <= 16'hFFFF;
rommem[11174] <= 16'hFFFF;
rommem[11175] <= 16'hFFFF;
rommem[11176] <= 16'hFFFF;
rommem[11177] <= 16'hFFFF;
rommem[11178] <= 16'hFFFF;
rommem[11179] <= 16'hFFFF;
rommem[11180] <= 16'hFFFF;
rommem[11181] <= 16'hFFFF;
rommem[11182] <= 16'hFFFF;
rommem[11183] <= 16'hFFFF;
rommem[11184] <= 16'hFFFF;
rommem[11185] <= 16'hFFFF;
rommem[11186] <= 16'hFFFF;
rommem[11187] <= 16'hFFFF;
rommem[11188] <= 16'hFFFF;
rommem[11189] <= 16'hFFFF;
rommem[11190] <= 16'hFFFF;
rommem[11191] <= 16'hFFFF;
rommem[11192] <= 16'hFFFF;
rommem[11193] <= 16'hFFFF;
rommem[11194] <= 16'hFFFF;
rommem[11195] <= 16'hFFFF;
rommem[11196] <= 16'hFFFF;
rommem[11197] <= 16'hFFFF;
rommem[11198] <= 16'hFFFF;
rommem[11199] <= 16'hFFFF;
rommem[11200] <= 16'hFFFF;
rommem[11201] <= 16'hFFFF;
rommem[11202] <= 16'hFFFF;
rommem[11203] <= 16'hFFFF;
rommem[11204] <= 16'hFFFF;
rommem[11205] <= 16'hFFFF;
rommem[11206] <= 16'hFFFF;
rommem[11207] <= 16'hFFFF;
rommem[11208] <= 16'hFFFF;
rommem[11209] <= 16'hFFFF;
rommem[11210] <= 16'hFFFF;
rommem[11211] <= 16'hFFFF;
rommem[11212] <= 16'hFFFF;
rommem[11213] <= 16'hFFFF;
rommem[11214] <= 16'hFFFF;
rommem[11215] <= 16'hFFFF;
rommem[11216] <= 16'hFFFF;
rommem[11217] <= 16'hFFFF;
rommem[11218] <= 16'hFFFF;
rommem[11219] <= 16'hFFFF;
rommem[11220] <= 16'hFFFF;
rommem[11221] <= 16'hFFFF;
rommem[11222] <= 16'hFFFF;
rommem[11223] <= 16'hFFFF;
rommem[11224] <= 16'hFFFF;
rommem[11225] <= 16'hFFFF;
rommem[11226] <= 16'hFFFF;
rommem[11227] <= 16'hFFFF;
rommem[11228] <= 16'hFFFF;
rommem[11229] <= 16'hFFFF;
rommem[11230] <= 16'hFFFF;
rommem[11231] <= 16'hFFFF;
rommem[11232] <= 16'hFFFF;
rommem[11233] <= 16'hFFFF;
rommem[11234] <= 16'hFFFF;
rommem[11235] <= 16'hFFFF;
rommem[11236] <= 16'hFFFF;
rommem[11237] <= 16'hFFFF;
rommem[11238] <= 16'hFFFF;
rommem[11239] <= 16'hFFFF;
rommem[11240] <= 16'hFFFF;
rommem[11241] <= 16'hFFFF;
rommem[11242] <= 16'hFFFF;
rommem[11243] <= 16'hFFFF;
rommem[11244] <= 16'hFFFF;
rommem[11245] <= 16'hFFFF;
rommem[11246] <= 16'hFFFF;
rommem[11247] <= 16'hFFFF;
rommem[11248] <= 16'hFFFF;
rommem[11249] <= 16'hFFFF;
rommem[11250] <= 16'hFFFF;
rommem[11251] <= 16'hFFFF;
rommem[11252] <= 16'hFFFF;
rommem[11253] <= 16'hFFFF;
rommem[11254] <= 16'hFFFF;
rommem[11255] <= 16'hFFFF;
rommem[11256] <= 16'hFFFF;
rommem[11257] <= 16'hFFFF;
rommem[11258] <= 16'hFFFF;
rommem[11259] <= 16'hFFFF;
rommem[11260] <= 16'hFFFF;
rommem[11261] <= 16'hFFFF;
rommem[11262] <= 16'hFFFF;
rommem[11263] <= 16'hFFFF;
rommem[11264] <= 16'hFFFF;
rommem[11265] <= 16'hFFFF;
rommem[11266] <= 16'hFFFF;
rommem[11267] <= 16'hFFFF;
rommem[11268] <= 16'hFFFF;
rommem[11269] <= 16'hFFFF;
rommem[11270] <= 16'hFFFF;
rommem[11271] <= 16'hFFFF;
rommem[11272] <= 16'hFFFF;
rommem[11273] <= 16'hFFFF;
rommem[11274] <= 16'hFFFF;
rommem[11275] <= 16'hFFFF;
rommem[11276] <= 16'hFFFF;
rommem[11277] <= 16'hFFFF;
rommem[11278] <= 16'hFFFF;
rommem[11279] <= 16'hFFFF;
rommem[11280] <= 16'hFFFF;
rommem[11281] <= 16'hFFFF;
rommem[11282] <= 16'hFFFF;
rommem[11283] <= 16'hFFFF;
rommem[11284] <= 16'hFFFF;
rommem[11285] <= 16'hFFFF;
rommem[11286] <= 16'hFFFF;
rommem[11287] <= 16'hFFFF;
rommem[11288] <= 16'hFFFF;
rommem[11289] <= 16'hFFFF;
rommem[11290] <= 16'hFFFF;
rommem[11291] <= 16'hFFFF;
rommem[11292] <= 16'hFFFF;
rommem[11293] <= 16'hFFFF;
rommem[11294] <= 16'hFFFF;
rommem[11295] <= 16'hFFFF;
rommem[11296] <= 16'hFFFF;
rommem[11297] <= 16'hFFFF;
rommem[11298] <= 16'hFFFF;
rommem[11299] <= 16'hFFFF;
rommem[11300] <= 16'hFFFF;
rommem[11301] <= 16'hFFFF;
rommem[11302] <= 16'hFFFF;
rommem[11303] <= 16'hFFFF;
rommem[11304] <= 16'hFFFF;
rommem[11305] <= 16'hFFFF;
rommem[11306] <= 16'hFFFF;
rommem[11307] <= 16'hFFFF;
rommem[11308] <= 16'hFFFF;
rommem[11309] <= 16'hFFFF;
rommem[11310] <= 16'hFFFF;
rommem[11311] <= 16'hFFFF;
rommem[11312] <= 16'hFFFF;
rommem[11313] <= 16'hFFFF;
rommem[11314] <= 16'hFFFF;
rommem[11315] <= 16'hFFFF;
rommem[11316] <= 16'hFFFF;
rommem[11317] <= 16'hFFFF;
rommem[11318] <= 16'hFFFF;
rommem[11319] <= 16'hFFFF;
rommem[11320] <= 16'hFFFF;
rommem[11321] <= 16'hFFFF;
rommem[11322] <= 16'hFFFF;
rommem[11323] <= 16'hFFFF;
rommem[11324] <= 16'hFFFF;
rommem[11325] <= 16'hFFFF;
rommem[11326] <= 16'hFFFF;
rommem[11327] <= 16'hFFFF;
rommem[11328] <= 16'hFFFF;
rommem[11329] <= 16'hFFFF;
rommem[11330] <= 16'hFFFF;
rommem[11331] <= 16'hFFFF;
rommem[11332] <= 16'hFFFF;
rommem[11333] <= 16'hFFFF;
rommem[11334] <= 16'hFFFF;
rommem[11335] <= 16'hFFFF;
rommem[11336] <= 16'hFFFF;
rommem[11337] <= 16'hFFFF;
rommem[11338] <= 16'hFFFF;
rommem[11339] <= 16'hFFFF;
rommem[11340] <= 16'hFFFF;
rommem[11341] <= 16'hFFFF;
rommem[11342] <= 16'hFFFF;
rommem[11343] <= 16'hFFFF;
rommem[11344] <= 16'hFFFF;
rommem[11345] <= 16'hFFFF;
rommem[11346] <= 16'hFFFF;
rommem[11347] <= 16'hFFFF;
rommem[11348] <= 16'hFFFF;
rommem[11349] <= 16'hFFFF;
rommem[11350] <= 16'hFFFF;
rommem[11351] <= 16'hFFFF;
rommem[11352] <= 16'hFFFF;
rommem[11353] <= 16'hFFFF;
rommem[11354] <= 16'hFFFF;
rommem[11355] <= 16'hFFFF;
rommem[11356] <= 16'hFFFF;
rommem[11357] <= 16'hFFFF;
rommem[11358] <= 16'hFFFF;
rommem[11359] <= 16'hFFFF;
rommem[11360] <= 16'hFFFF;
rommem[11361] <= 16'hFFFF;
rommem[11362] <= 16'hFFFF;
rommem[11363] <= 16'hFFFF;
rommem[11364] <= 16'hFFFF;
rommem[11365] <= 16'hFFFF;
rommem[11366] <= 16'hFFFF;
rommem[11367] <= 16'hFFFF;
rommem[11368] <= 16'hFFFF;
rommem[11369] <= 16'hFFFF;
rommem[11370] <= 16'hFFFF;
rommem[11371] <= 16'hFFFF;
rommem[11372] <= 16'hFFFF;
rommem[11373] <= 16'hFFFF;
rommem[11374] <= 16'hFFFF;
rommem[11375] <= 16'hFFFF;
rommem[11376] <= 16'hFFFF;
rommem[11377] <= 16'hFFFF;
rommem[11378] <= 16'hFFFF;
rommem[11379] <= 16'hFFFF;
rommem[11380] <= 16'hFFFF;
rommem[11381] <= 16'hFFFF;
rommem[11382] <= 16'hFFFF;
rommem[11383] <= 16'hFFFF;
rommem[11384] <= 16'hFFFF;
rommem[11385] <= 16'hFFFF;
rommem[11386] <= 16'hFFFF;
rommem[11387] <= 16'hFFFF;
rommem[11388] <= 16'hFFFF;
rommem[11389] <= 16'hFFFF;
rommem[11390] <= 16'hFFFF;
rommem[11391] <= 16'hFFFF;
rommem[11392] <= 16'hFFFF;
rommem[11393] <= 16'hFFFF;
rommem[11394] <= 16'hFFFF;
rommem[11395] <= 16'hFFFF;
rommem[11396] <= 16'hFFFF;
rommem[11397] <= 16'hFFFF;
rommem[11398] <= 16'hFFFF;
rommem[11399] <= 16'hFFFF;
rommem[11400] <= 16'hFFFF;
rommem[11401] <= 16'hFFFF;
rommem[11402] <= 16'hFFFF;
rommem[11403] <= 16'hFFFF;
rommem[11404] <= 16'hFFFF;
rommem[11405] <= 16'hFFFF;
rommem[11406] <= 16'hFFFF;
rommem[11407] <= 16'hFFFF;
rommem[11408] <= 16'hFFFF;
rommem[11409] <= 16'hFFFF;
rommem[11410] <= 16'hFFFF;
rommem[11411] <= 16'hFFFF;
rommem[11412] <= 16'hFFFF;
rommem[11413] <= 16'hFFFF;
rommem[11414] <= 16'hFFFF;
rommem[11415] <= 16'hFFFF;
rommem[11416] <= 16'hFFFF;
rommem[11417] <= 16'hFFFF;
rommem[11418] <= 16'hFFFF;
rommem[11419] <= 16'hFFFF;
rommem[11420] <= 16'hFFFF;
rommem[11421] <= 16'hFFFF;
rommem[11422] <= 16'hFFFF;
rommem[11423] <= 16'hFFFF;
rommem[11424] <= 16'hFFFF;
rommem[11425] <= 16'hFFFF;
rommem[11426] <= 16'hFFFF;
rommem[11427] <= 16'hFFFF;
rommem[11428] <= 16'hFFFF;
rommem[11429] <= 16'hFFFF;
rommem[11430] <= 16'hFFFF;
rommem[11431] <= 16'hFFFF;
rommem[11432] <= 16'hFFFF;
rommem[11433] <= 16'hFFFF;
rommem[11434] <= 16'hFFFF;
rommem[11435] <= 16'hFFFF;
rommem[11436] <= 16'hFFFF;
rommem[11437] <= 16'hFFFF;
rommem[11438] <= 16'hFFFF;
rommem[11439] <= 16'hFFFF;
rommem[11440] <= 16'hFFFF;
rommem[11441] <= 16'hFFFF;
rommem[11442] <= 16'hFFFF;
rommem[11443] <= 16'hFFFF;
rommem[11444] <= 16'hFFFF;
rommem[11445] <= 16'hFFFF;
rommem[11446] <= 16'hFFFF;
rommem[11447] <= 16'hFFFF;
rommem[11448] <= 16'hFFFF;
rommem[11449] <= 16'hFFFF;
rommem[11450] <= 16'hFFFF;
rommem[11451] <= 16'hFFFF;
rommem[11452] <= 16'hFFFF;
rommem[11453] <= 16'hFFFF;
rommem[11454] <= 16'hFFFF;
rommem[11455] <= 16'hFFFF;
rommem[11456] <= 16'hFFFF;
rommem[11457] <= 16'hFFFF;
rommem[11458] <= 16'hFFFF;
rommem[11459] <= 16'hFFFF;
rommem[11460] <= 16'hFFFF;
rommem[11461] <= 16'hFFFF;
rommem[11462] <= 16'hFFFF;
rommem[11463] <= 16'hFFFF;
rommem[11464] <= 16'hFFFF;
rommem[11465] <= 16'hFFFF;
rommem[11466] <= 16'hFFFF;
rommem[11467] <= 16'hFFFF;
rommem[11468] <= 16'hFFFF;
rommem[11469] <= 16'hFFFF;
rommem[11470] <= 16'hFFFF;
rommem[11471] <= 16'hFFFF;
rommem[11472] <= 16'hFFFF;
rommem[11473] <= 16'hFFFF;
rommem[11474] <= 16'hFFFF;
rommem[11475] <= 16'hFFFF;
rommem[11476] <= 16'hFFFF;
rommem[11477] <= 16'hFFFF;
rommem[11478] <= 16'hFFFF;
rommem[11479] <= 16'hFFFF;
rommem[11480] <= 16'hFFFF;
rommem[11481] <= 16'hFFFF;
rommem[11482] <= 16'hFFFF;
rommem[11483] <= 16'hFFFF;
rommem[11484] <= 16'hFFFF;
rommem[11485] <= 16'hFFFF;
rommem[11486] <= 16'hFFFF;
rommem[11487] <= 16'hFFFF;
rommem[11488] <= 16'hFFFF;
rommem[11489] <= 16'hFFFF;
rommem[11490] <= 16'hFFFF;
rommem[11491] <= 16'hFFFF;
rommem[11492] <= 16'hFFFF;
rommem[11493] <= 16'hFFFF;
rommem[11494] <= 16'hFFFF;
rommem[11495] <= 16'hFFFF;
rommem[11496] <= 16'hFFFF;
rommem[11497] <= 16'hFFFF;
rommem[11498] <= 16'hFFFF;
rommem[11499] <= 16'hFFFF;
rommem[11500] <= 16'hFFFF;
rommem[11501] <= 16'hFFFF;
rommem[11502] <= 16'hFFFF;
rommem[11503] <= 16'hFFFF;
rommem[11504] <= 16'hFFFF;
rommem[11505] <= 16'hFFFF;
rommem[11506] <= 16'hFFFF;
rommem[11507] <= 16'hFFFF;
rommem[11508] <= 16'hFFFF;
rommem[11509] <= 16'hFFFF;
rommem[11510] <= 16'hFFFF;
rommem[11511] <= 16'hFFFF;
rommem[11512] <= 16'hFFFF;
rommem[11513] <= 16'hFFFF;
rommem[11514] <= 16'hFFFF;
rommem[11515] <= 16'hFFFF;
rommem[11516] <= 16'hFFFF;
rommem[11517] <= 16'hFFFF;
rommem[11518] <= 16'hFFFF;
rommem[11519] <= 16'hFFFF;
rommem[11520] <= 16'hFFFF;
rommem[11521] <= 16'hFFFF;
rommem[11522] <= 16'hFFFF;
rommem[11523] <= 16'hFFFF;
rommem[11524] <= 16'hFFFF;
rommem[11525] <= 16'hFFFF;
rommem[11526] <= 16'hFFFF;
rommem[11527] <= 16'hFFFF;
rommem[11528] <= 16'hFFFF;
rommem[11529] <= 16'hFFFF;
rommem[11530] <= 16'hFFFF;
rommem[11531] <= 16'hFFFF;
rommem[11532] <= 16'hFFFF;
rommem[11533] <= 16'hFFFF;
rommem[11534] <= 16'hFFFF;
rommem[11535] <= 16'hFFFF;
rommem[11536] <= 16'hFFFF;
rommem[11537] <= 16'hFFFF;
rommem[11538] <= 16'hFFFF;
rommem[11539] <= 16'hFFFF;
rommem[11540] <= 16'hFFFF;
rommem[11541] <= 16'hFFFF;
rommem[11542] <= 16'hFFFF;
rommem[11543] <= 16'hFFFF;
rommem[11544] <= 16'hFFFF;
rommem[11545] <= 16'hFFFF;
rommem[11546] <= 16'hFFFF;
rommem[11547] <= 16'hFFFF;
rommem[11548] <= 16'hFFFF;
rommem[11549] <= 16'hFFFF;
rommem[11550] <= 16'hFFFF;
rommem[11551] <= 16'hFFFF;
rommem[11552] <= 16'hFFFF;
rommem[11553] <= 16'hFFFF;
rommem[11554] <= 16'hFFFF;
rommem[11555] <= 16'hFFFF;
rommem[11556] <= 16'hFFFF;
rommem[11557] <= 16'hFFFF;
rommem[11558] <= 16'hFFFF;
rommem[11559] <= 16'hFFFF;
rommem[11560] <= 16'hFFFF;
rommem[11561] <= 16'hFFFF;
rommem[11562] <= 16'hFFFF;
rommem[11563] <= 16'hFFFF;
rommem[11564] <= 16'hFFFF;
rommem[11565] <= 16'hFFFF;
rommem[11566] <= 16'hFFFF;
rommem[11567] <= 16'hFFFF;
rommem[11568] <= 16'hFFFF;
rommem[11569] <= 16'hFFFF;
rommem[11570] <= 16'hFFFF;
rommem[11571] <= 16'hFFFF;
rommem[11572] <= 16'hFFFF;
rommem[11573] <= 16'hFFFF;
rommem[11574] <= 16'hFFFF;
rommem[11575] <= 16'hFFFF;
rommem[11576] <= 16'hFFFF;
rommem[11577] <= 16'hFFFF;
rommem[11578] <= 16'hFFFF;
rommem[11579] <= 16'hFFFF;
rommem[11580] <= 16'hFFFF;
rommem[11581] <= 16'hFFFF;
rommem[11582] <= 16'hFFFF;
rommem[11583] <= 16'hFFFF;
rommem[11584] <= 16'hFFFF;
rommem[11585] <= 16'hFFFF;
rommem[11586] <= 16'hFFFF;
rommem[11587] <= 16'hFFFF;
rommem[11588] <= 16'hFFFF;
rommem[11589] <= 16'hFFFF;
rommem[11590] <= 16'hFFFF;
rommem[11591] <= 16'hFFFF;
rommem[11592] <= 16'hFFFF;
rommem[11593] <= 16'hFFFF;
rommem[11594] <= 16'hFFFF;
rommem[11595] <= 16'hFFFF;
rommem[11596] <= 16'hFFFF;
rommem[11597] <= 16'hFFFF;
rommem[11598] <= 16'hFFFF;
rommem[11599] <= 16'hFFFF;
rommem[11600] <= 16'hFFFF;
rommem[11601] <= 16'hFFFF;
rommem[11602] <= 16'hFFFF;
rommem[11603] <= 16'hFFFF;
rommem[11604] <= 16'hFFFF;
rommem[11605] <= 16'hFFFF;
rommem[11606] <= 16'hFFFF;
rommem[11607] <= 16'hFFFF;
rommem[11608] <= 16'hFFFF;
rommem[11609] <= 16'hFFFF;
rommem[11610] <= 16'hFFFF;
rommem[11611] <= 16'hFFFF;
rommem[11612] <= 16'hFFFF;
rommem[11613] <= 16'hFFFF;
rommem[11614] <= 16'hFFFF;
rommem[11615] <= 16'hFFFF;
rommem[11616] <= 16'hFFFF;
rommem[11617] <= 16'hFFFF;
rommem[11618] <= 16'hFFFF;
rommem[11619] <= 16'hFFFF;
rommem[11620] <= 16'hFFFF;
rommem[11621] <= 16'hFFFF;
rommem[11622] <= 16'hFFFF;
rommem[11623] <= 16'hFFFF;
rommem[11624] <= 16'hFFFF;
rommem[11625] <= 16'hFFFF;
rommem[11626] <= 16'hFFFF;
rommem[11627] <= 16'hFFFF;
rommem[11628] <= 16'hFFFF;
rommem[11629] <= 16'hFFFF;
rommem[11630] <= 16'hFFFF;
rommem[11631] <= 16'hFFFF;
rommem[11632] <= 16'hFFFF;
rommem[11633] <= 16'hFFFF;
rommem[11634] <= 16'hFFFF;
rommem[11635] <= 16'hFFFF;
rommem[11636] <= 16'hFFFF;
rommem[11637] <= 16'hFFFF;
rommem[11638] <= 16'hFFFF;
rommem[11639] <= 16'hFFFF;
rommem[11640] <= 16'hFFFF;
rommem[11641] <= 16'hFFFF;
rommem[11642] <= 16'hFFFF;
rommem[11643] <= 16'hFFFF;
rommem[11644] <= 16'hFFFF;
rommem[11645] <= 16'hFFFF;
rommem[11646] <= 16'hFFFF;
rommem[11647] <= 16'hFFFF;
rommem[11648] <= 16'hFFFF;
rommem[11649] <= 16'hFFFF;
rommem[11650] <= 16'hFFFF;
rommem[11651] <= 16'hFFFF;
rommem[11652] <= 16'hFFFF;
rommem[11653] <= 16'hFFFF;
rommem[11654] <= 16'hFFFF;
rommem[11655] <= 16'hFFFF;
rommem[11656] <= 16'hFFFF;
rommem[11657] <= 16'hFFFF;
rommem[11658] <= 16'hFFFF;
rommem[11659] <= 16'hFFFF;
rommem[11660] <= 16'hFFFF;
rommem[11661] <= 16'hFFFF;
rommem[11662] <= 16'hFFFF;
rommem[11663] <= 16'hFFFF;
rommem[11664] <= 16'hFFFF;
rommem[11665] <= 16'hFFFF;
rommem[11666] <= 16'hFFFF;
rommem[11667] <= 16'hFFFF;
rommem[11668] <= 16'hFFFF;
rommem[11669] <= 16'hFFFF;
rommem[11670] <= 16'hFFFF;
rommem[11671] <= 16'hFFFF;
rommem[11672] <= 16'hFFFF;
rommem[11673] <= 16'hFFFF;
rommem[11674] <= 16'hFFFF;
rommem[11675] <= 16'hFFFF;
rommem[11676] <= 16'hFFFF;
rommem[11677] <= 16'hFFFF;
rommem[11678] <= 16'hFFFF;
rommem[11679] <= 16'hFFFF;
rommem[11680] <= 16'hFFFF;
rommem[11681] <= 16'hFFFF;
rommem[11682] <= 16'hFFFF;
rommem[11683] <= 16'hFFFF;
rommem[11684] <= 16'hFFFF;
rommem[11685] <= 16'hFFFF;
rommem[11686] <= 16'hFFFF;
rommem[11687] <= 16'hFFFF;
rommem[11688] <= 16'hFFFF;
rommem[11689] <= 16'hFFFF;
rommem[11690] <= 16'hFFFF;
rommem[11691] <= 16'hFFFF;
rommem[11692] <= 16'hFFFF;
rommem[11693] <= 16'hFFFF;
rommem[11694] <= 16'hFFFF;
rommem[11695] <= 16'hFFFF;
rommem[11696] <= 16'hFFFF;
rommem[11697] <= 16'hFFFF;
rommem[11698] <= 16'hFFFF;
rommem[11699] <= 16'hFFFF;
rommem[11700] <= 16'hFFFF;
rommem[11701] <= 16'hFFFF;
rommem[11702] <= 16'hFFFF;
rommem[11703] <= 16'hFFFF;
rommem[11704] <= 16'hFFFF;
rommem[11705] <= 16'hFFFF;
rommem[11706] <= 16'hFFFF;
rommem[11707] <= 16'hFFFF;
rommem[11708] <= 16'hFFFF;
rommem[11709] <= 16'hFFFF;
rommem[11710] <= 16'hFFFF;
rommem[11711] <= 16'hFFFF;
rommem[11712] <= 16'hFFFF;
rommem[11713] <= 16'hFFFF;
rommem[11714] <= 16'hFFFF;
rommem[11715] <= 16'hFFFF;
rommem[11716] <= 16'hFFFF;
rommem[11717] <= 16'hFFFF;
rommem[11718] <= 16'hFFFF;
rommem[11719] <= 16'hFFFF;
rommem[11720] <= 16'hFFFF;
rommem[11721] <= 16'hFFFF;
rommem[11722] <= 16'hFFFF;
rommem[11723] <= 16'hFFFF;
rommem[11724] <= 16'hFFFF;
rommem[11725] <= 16'hFFFF;
rommem[11726] <= 16'hFFFF;
rommem[11727] <= 16'hFFFF;
rommem[11728] <= 16'hFFFF;
rommem[11729] <= 16'hFFFF;
rommem[11730] <= 16'hFFFF;
rommem[11731] <= 16'hFFFF;
rommem[11732] <= 16'hFFFF;
rommem[11733] <= 16'hFFFF;
rommem[11734] <= 16'hFFFF;
rommem[11735] <= 16'hFFFF;
rommem[11736] <= 16'hFFFF;
rommem[11737] <= 16'hFFFF;
rommem[11738] <= 16'hFFFF;
rommem[11739] <= 16'hFFFF;
rommem[11740] <= 16'hFFFF;
rommem[11741] <= 16'hFFFF;
rommem[11742] <= 16'hFFFF;
rommem[11743] <= 16'hFFFF;
rommem[11744] <= 16'hFFFF;
rommem[11745] <= 16'hFFFF;
rommem[11746] <= 16'hFFFF;
rommem[11747] <= 16'hFFFF;
rommem[11748] <= 16'hFFFF;
rommem[11749] <= 16'hFFFF;
rommem[11750] <= 16'hFFFF;
rommem[11751] <= 16'hFFFF;
rommem[11752] <= 16'hFFFF;
rommem[11753] <= 16'hFFFF;
rommem[11754] <= 16'hFFFF;
rommem[11755] <= 16'hFFFF;
rommem[11756] <= 16'hFFFF;
rommem[11757] <= 16'hFFFF;
rommem[11758] <= 16'hFFFF;
rommem[11759] <= 16'hFFFF;
rommem[11760] <= 16'hFFFF;
rommem[11761] <= 16'hFFFF;
rommem[11762] <= 16'hFFFF;
rommem[11763] <= 16'hFFFF;
rommem[11764] <= 16'hFFFF;
rommem[11765] <= 16'hFFFF;
rommem[11766] <= 16'hFFFF;
rommem[11767] <= 16'hFFFF;
rommem[11768] <= 16'hFFFF;
rommem[11769] <= 16'hFFFF;
rommem[11770] <= 16'hFFFF;
rommem[11771] <= 16'hFFFF;
rommem[11772] <= 16'hFFFF;
rommem[11773] <= 16'hFFFF;
rommem[11774] <= 16'hFFFF;
rommem[11775] <= 16'hFFFF;
rommem[11776] <= 16'hFFFF;
rommem[11777] <= 16'hFFFF;
rommem[11778] <= 16'hFFFF;
rommem[11779] <= 16'hFFFF;
rommem[11780] <= 16'hFFFF;
rommem[11781] <= 16'hFFFF;
rommem[11782] <= 16'hFFFF;
rommem[11783] <= 16'hFFFF;
rommem[11784] <= 16'hFFFF;
rommem[11785] <= 16'hFFFF;
rommem[11786] <= 16'hFFFF;
rommem[11787] <= 16'hFFFF;
rommem[11788] <= 16'hFFFF;
rommem[11789] <= 16'hFFFF;
rommem[11790] <= 16'hFFFF;
rommem[11791] <= 16'hFFFF;
rommem[11792] <= 16'hFFFF;
rommem[11793] <= 16'hFFFF;
rommem[11794] <= 16'hFFFF;
rommem[11795] <= 16'hFFFF;
rommem[11796] <= 16'hFFFF;
rommem[11797] <= 16'hFFFF;
rommem[11798] <= 16'hFFFF;
rommem[11799] <= 16'hFFFF;
rommem[11800] <= 16'hFFFF;
rommem[11801] <= 16'hFFFF;
rommem[11802] <= 16'hFFFF;
rommem[11803] <= 16'hFFFF;
rommem[11804] <= 16'hFFFF;
rommem[11805] <= 16'hFFFF;
rommem[11806] <= 16'hFFFF;
rommem[11807] <= 16'hFFFF;
rommem[11808] <= 16'hFFFF;
rommem[11809] <= 16'hFFFF;
rommem[11810] <= 16'hFFFF;
rommem[11811] <= 16'hFFFF;
rommem[11812] <= 16'hFFFF;
rommem[11813] <= 16'hFFFF;
rommem[11814] <= 16'hFFFF;
rommem[11815] <= 16'hFFFF;
rommem[11816] <= 16'hFFFF;
rommem[11817] <= 16'hFFFF;
rommem[11818] <= 16'hFFFF;
rommem[11819] <= 16'hFFFF;
rommem[11820] <= 16'hFFFF;
rommem[11821] <= 16'hFFFF;
rommem[11822] <= 16'hFFFF;
rommem[11823] <= 16'hFFFF;
rommem[11824] <= 16'hFFFF;
rommem[11825] <= 16'hFFFF;
rommem[11826] <= 16'hFFFF;
rommem[11827] <= 16'hFFFF;
rommem[11828] <= 16'hFFFF;
rommem[11829] <= 16'hFFFF;
rommem[11830] <= 16'hFFFF;
rommem[11831] <= 16'hFFFF;
rommem[11832] <= 16'hFFFF;
rommem[11833] <= 16'hFFFF;
rommem[11834] <= 16'hFFFF;
rommem[11835] <= 16'hFFFF;
rommem[11836] <= 16'hFFFF;
rommem[11837] <= 16'hFFFF;
rommem[11838] <= 16'hFFFF;
rommem[11839] <= 16'hFFFF;
rommem[11840] <= 16'hFFFF;
rommem[11841] <= 16'hFFFF;
rommem[11842] <= 16'hFFFF;
rommem[11843] <= 16'hFFFF;
rommem[11844] <= 16'hFFFF;
rommem[11845] <= 16'hFFFF;
rommem[11846] <= 16'hFFFF;
rommem[11847] <= 16'hFFFF;
rommem[11848] <= 16'hFFFF;
rommem[11849] <= 16'hFFFF;
rommem[11850] <= 16'hFFFF;
rommem[11851] <= 16'hFFFF;
rommem[11852] <= 16'hFFFF;
rommem[11853] <= 16'hFFFF;
rommem[11854] <= 16'hFFFF;
rommem[11855] <= 16'hFFFF;
rommem[11856] <= 16'hFFFF;
rommem[11857] <= 16'hFFFF;
rommem[11858] <= 16'hFFFF;
rommem[11859] <= 16'hFFFF;
rommem[11860] <= 16'hFFFF;
rommem[11861] <= 16'hFFFF;
rommem[11862] <= 16'hFFFF;
rommem[11863] <= 16'hFFFF;
rommem[11864] <= 16'hFFFF;
rommem[11865] <= 16'hFFFF;
rommem[11866] <= 16'hFFFF;
rommem[11867] <= 16'hFFFF;
rommem[11868] <= 16'hFFFF;
rommem[11869] <= 16'hFFFF;
rommem[11870] <= 16'hFFFF;
rommem[11871] <= 16'hFFFF;
rommem[11872] <= 16'hFFFF;
rommem[11873] <= 16'hFFFF;
rommem[11874] <= 16'hFFFF;
rommem[11875] <= 16'hFFFF;
rommem[11876] <= 16'hFFFF;
rommem[11877] <= 16'hFFFF;
rommem[11878] <= 16'hFFFF;
rommem[11879] <= 16'hFFFF;
rommem[11880] <= 16'hFFFF;
rommem[11881] <= 16'hFFFF;
rommem[11882] <= 16'hFFFF;
rommem[11883] <= 16'hFFFF;
rommem[11884] <= 16'hFFFF;
rommem[11885] <= 16'hFFFF;
rommem[11886] <= 16'hFFFF;
rommem[11887] <= 16'hFFFF;
rommem[11888] <= 16'hFFFF;
rommem[11889] <= 16'hFFFF;
rommem[11890] <= 16'hFFFF;
rommem[11891] <= 16'hFFFF;
rommem[11892] <= 16'hFFFF;
rommem[11893] <= 16'hFFFF;
rommem[11894] <= 16'hFFFF;
rommem[11895] <= 16'hFFFF;
rommem[11896] <= 16'hFFFF;
rommem[11897] <= 16'hFFFF;
rommem[11898] <= 16'hFFFF;
rommem[11899] <= 16'hFFFF;
rommem[11900] <= 16'hFFFF;
rommem[11901] <= 16'hFFFF;
rommem[11902] <= 16'hFFFF;
rommem[11903] <= 16'hFFFF;
rommem[11904] <= 16'hFFFF;
rommem[11905] <= 16'hFFFF;
rommem[11906] <= 16'hFFFF;
rommem[11907] <= 16'hFFFF;
rommem[11908] <= 16'hFFFF;
rommem[11909] <= 16'hFFFF;
rommem[11910] <= 16'hFFFF;
rommem[11911] <= 16'hFFFF;
rommem[11912] <= 16'hFFFF;
rommem[11913] <= 16'hFFFF;
rommem[11914] <= 16'hFFFF;
rommem[11915] <= 16'hFFFF;
rommem[11916] <= 16'hFFFF;
rommem[11917] <= 16'hFFFF;
rommem[11918] <= 16'hFFFF;
rommem[11919] <= 16'hFFFF;
rommem[11920] <= 16'hFFFF;
rommem[11921] <= 16'hFFFF;
rommem[11922] <= 16'hFFFF;
rommem[11923] <= 16'hFFFF;
rommem[11924] <= 16'hFFFF;
rommem[11925] <= 16'hFFFF;
rommem[11926] <= 16'hFFFF;
rommem[11927] <= 16'hFFFF;
rommem[11928] <= 16'hFFFF;
rommem[11929] <= 16'hFFFF;
rommem[11930] <= 16'hFFFF;
rommem[11931] <= 16'hFFFF;
rommem[11932] <= 16'hFFFF;
rommem[11933] <= 16'hFFFF;
rommem[11934] <= 16'hFFFF;
rommem[11935] <= 16'hFFFF;
rommem[11936] <= 16'hFFFF;
rommem[11937] <= 16'hFFFF;
rommem[11938] <= 16'hFFFF;
rommem[11939] <= 16'hFFFF;
rommem[11940] <= 16'hFFFF;
rommem[11941] <= 16'hFFFF;
rommem[11942] <= 16'hFFFF;
rommem[11943] <= 16'hFFFF;
rommem[11944] <= 16'hFFFF;
rommem[11945] <= 16'hFFFF;
rommem[11946] <= 16'hFFFF;
rommem[11947] <= 16'hFFFF;
rommem[11948] <= 16'hFFFF;
rommem[11949] <= 16'hFFFF;
rommem[11950] <= 16'hFFFF;
rommem[11951] <= 16'hFFFF;
rommem[11952] <= 16'hFFFF;
rommem[11953] <= 16'hFFFF;
rommem[11954] <= 16'hFFFF;
rommem[11955] <= 16'hFFFF;
rommem[11956] <= 16'hFFFF;
rommem[11957] <= 16'hFFFF;
rommem[11958] <= 16'hFFFF;
rommem[11959] <= 16'hFFFF;
rommem[11960] <= 16'hFFFF;
rommem[11961] <= 16'hFFFF;
rommem[11962] <= 16'hFFFF;
rommem[11963] <= 16'hFFFF;
rommem[11964] <= 16'hFFFF;
rommem[11965] <= 16'hFFFF;
rommem[11966] <= 16'hFFFF;
rommem[11967] <= 16'hFFFF;
rommem[11968] <= 16'hFFFF;
rommem[11969] <= 16'hFFFF;
rommem[11970] <= 16'hFFFF;
rommem[11971] <= 16'hFFFF;
rommem[11972] <= 16'hFFFF;
rommem[11973] <= 16'hFFFF;
rommem[11974] <= 16'hFFFF;
rommem[11975] <= 16'hFFFF;
rommem[11976] <= 16'hFFFF;
rommem[11977] <= 16'hFFFF;
rommem[11978] <= 16'hFFFF;
rommem[11979] <= 16'hFFFF;
rommem[11980] <= 16'hFFFF;
rommem[11981] <= 16'hFFFF;
rommem[11982] <= 16'hFFFF;
rommem[11983] <= 16'hFFFF;
rommem[11984] <= 16'hFFFF;
rommem[11985] <= 16'hFFFF;
rommem[11986] <= 16'hFFFF;
rommem[11987] <= 16'hFFFF;
rommem[11988] <= 16'hFFFF;
rommem[11989] <= 16'hFFFF;
rommem[11990] <= 16'hFFFF;
rommem[11991] <= 16'hFFFF;
rommem[11992] <= 16'hFFFF;
rommem[11993] <= 16'hFFFF;
rommem[11994] <= 16'hFFFF;
rommem[11995] <= 16'hFFFF;
rommem[11996] <= 16'hFFFF;
rommem[11997] <= 16'hFFFF;
rommem[11998] <= 16'hFFFF;
rommem[11999] <= 16'hFFFF;
rommem[12000] <= 16'hFFFF;
rommem[12001] <= 16'hFFFF;
rommem[12002] <= 16'hFFFF;
rommem[12003] <= 16'hFFFF;
rommem[12004] <= 16'hFFFF;
rommem[12005] <= 16'hFFFF;
rommem[12006] <= 16'hFFFF;
rommem[12007] <= 16'hFFFF;
rommem[12008] <= 16'hFFFF;
rommem[12009] <= 16'hFFFF;
rommem[12010] <= 16'hFFFF;
rommem[12011] <= 16'hFFFF;
rommem[12012] <= 16'hFFFF;
rommem[12013] <= 16'hFFFF;
rommem[12014] <= 16'hFFFF;
rommem[12015] <= 16'hFFFF;
rommem[12016] <= 16'hFFFF;
rommem[12017] <= 16'hFFFF;
rommem[12018] <= 16'hFFFF;
rommem[12019] <= 16'hFFFF;
rommem[12020] <= 16'hFFFF;
rommem[12021] <= 16'hFFFF;
rommem[12022] <= 16'hFFFF;
rommem[12023] <= 16'hFFFF;
rommem[12024] <= 16'hFFFF;
rommem[12025] <= 16'hFFFF;
rommem[12026] <= 16'hFFFF;
rommem[12027] <= 16'hFFFF;
rommem[12028] <= 16'hFFFF;
rommem[12029] <= 16'hFFFF;
rommem[12030] <= 16'hFFFF;
rommem[12031] <= 16'hFFFF;
rommem[12032] <= 16'hFFFF;
rommem[12033] <= 16'hFFFF;
rommem[12034] <= 16'hFFFF;
rommem[12035] <= 16'hFFFF;
rommem[12036] <= 16'hFFFF;
rommem[12037] <= 16'hFFFF;
rommem[12038] <= 16'hFFFF;
rommem[12039] <= 16'hFFFF;
rommem[12040] <= 16'hFFFF;
rommem[12041] <= 16'hFFFF;
rommem[12042] <= 16'hFFFF;
rommem[12043] <= 16'hFFFF;
rommem[12044] <= 16'hFFFF;
rommem[12045] <= 16'hFFFF;
rommem[12046] <= 16'hFFFF;
rommem[12047] <= 16'hFFFF;
rommem[12048] <= 16'hFFFF;
rommem[12049] <= 16'hFFFF;
rommem[12050] <= 16'hFFFF;
rommem[12051] <= 16'hFFFF;
rommem[12052] <= 16'hFFFF;
rommem[12053] <= 16'hFFFF;
rommem[12054] <= 16'hFFFF;
rommem[12055] <= 16'hFFFF;
rommem[12056] <= 16'hFFFF;
rommem[12057] <= 16'hFFFF;
rommem[12058] <= 16'hFFFF;
rommem[12059] <= 16'hFFFF;
rommem[12060] <= 16'hFFFF;
rommem[12061] <= 16'hFFFF;
rommem[12062] <= 16'hFFFF;
rommem[12063] <= 16'hFFFF;
rommem[12064] <= 16'hFFFF;
rommem[12065] <= 16'hFFFF;
rommem[12066] <= 16'hFFFF;
rommem[12067] <= 16'hFFFF;
rommem[12068] <= 16'hFFFF;
rommem[12069] <= 16'hFFFF;
rommem[12070] <= 16'hFFFF;
rommem[12071] <= 16'hFFFF;
rommem[12072] <= 16'hFFFF;
rommem[12073] <= 16'hFFFF;
rommem[12074] <= 16'hFFFF;
rommem[12075] <= 16'hFFFF;
rommem[12076] <= 16'hFFFF;
rommem[12077] <= 16'hFFFF;
rommem[12078] <= 16'hFFFF;
rommem[12079] <= 16'hFFFF;
rommem[12080] <= 16'hFFFF;
rommem[12081] <= 16'hFFFF;
rommem[12082] <= 16'hFFFF;
rommem[12083] <= 16'hFFFF;
rommem[12084] <= 16'hFFFF;
rommem[12085] <= 16'hFFFF;
rommem[12086] <= 16'hFFFF;
rommem[12087] <= 16'hFFFF;
rommem[12088] <= 16'hFFFF;
rommem[12089] <= 16'hFFFF;
rommem[12090] <= 16'hFFFF;
rommem[12091] <= 16'hFFFF;
rommem[12092] <= 16'hFFFF;
rommem[12093] <= 16'hFFFF;
rommem[12094] <= 16'hFFFF;
rommem[12095] <= 16'hFFFF;
rommem[12096] <= 16'hFFFF;
rommem[12097] <= 16'hFFFF;
rommem[12098] <= 16'hFFFF;
rommem[12099] <= 16'hFFFF;
rommem[12100] <= 16'hFFFF;
rommem[12101] <= 16'hFFFF;
rommem[12102] <= 16'hFFFF;
rommem[12103] <= 16'hFFFF;
rommem[12104] <= 16'hFFFF;
rommem[12105] <= 16'hFFFF;
rommem[12106] <= 16'hFFFF;
rommem[12107] <= 16'hFFFF;
rommem[12108] <= 16'hFFFF;
rommem[12109] <= 16'hFFFF;
rommem[12110] <= 16'hFFFF;
rommem[12111] <= 16'hFFFF;
rommem[12112] <= 16'hFFFF;
rommem[12113] <= 16'hFFFF;
rommem[12114] <= 16'hFFFF;
rommem[12115] <= 16'hFFFF;
rommem[12116] <= 16'hFFFF;
rommem[12117] <= 16'hFFFF;
rommem[12118] <= 16'hFFFF;
rommem[12119] <= 16'hFFFF;
rommem[12120] <= 16'hFFFF;
rommem[12121] <= 16'hFFFF;
rommem[12122] <= 16'hFFFF;
rommem[12123] <= 16'hFFFF;
rommem[12124] <= 16'hFFFF;
rommem[12125] <= 16'hFFFF;
rommem[12126] <= 16'hFFFF;
rommem[12127] <= 16'hFFFF;
rommem[12128] <= 16'hFFFF;
rommem[12129] <= 16'hFFFF;
rommem[12130] <= 16'hFFFF;
rommem[12131] <= 16'hFFFF;
rommem[12132] <= 16'hFFFF;
rommem[12133] <= 16'hFFFF;
rommem[12134] <= 16'hFFFF;
rommem[12135] <= 16'hFFFF;
rommem[12136] <= 16'hFFFF;
rommem[12137] <= 16'hFFFF;
rommem[12138] <= 16'hFFFF;
rommem[12139] <= 16'hFFFF;
rommem[12140] <= 16'hFFFF;
rommem[12141] <= 16'hFFFF;
rommem[12142] <= 16'hFFFF;
rommem[12143] <= 16'hFFFF;
rommem[12144] <= 16'hFFFF;
rommem[12145] <= 16'hFFFF;
rommem[12146] <= 16'hFFFF;
rommem[12147] <= 16'hFFFF;
rommem[12148] <= 16'hFFFF;
rommem[12149] <= 16'hFFFF;
rommem[12150] <= 16'hFFFF;
rommem[12151] <= 16'hFFFF;
rommem[12152] <= 16'hFFFF;
rommem[12153] <= 16'hFFFF;
rommem[12154] <= 16'hFFFF;
rommem[12155] <= 16'hFFFF;
rommem[12156] <= 16'hFFFF;
rommem[12157] <= 16'hFFFF;
rommem[12158] <= 16'hFFFF;
rommem[12159] <= 16'hFFFF;
rommem[12160] <= 16'hFFFF;
rommem[12161] <= 16'hFFFF;
rommem[12162] <= 16'hFFFF;
rommem[12163] <= 16'hFFFF;
rommem[12164] <= 16'hFFFF;
rommem[12165] <= 16'hFFFF;
rommem[12166] <= 16'hFFFF;
rommem[12167] <= 16'hFFFF;
rommem[12168] <= 16'hFFFF;
rommem[12169] <= 16'hFFFF;
rommem[12170] <= 16'hFFFF;
rommem[12171] <= 16'hFFFF;
rommem[12172] <= 16'hFFFF;
rommem[12173] <= 16'hFFFF;
rommem[12174] <= 16'hFFFF;
rommem[12175] <= 16'hFFFF;
rommem[12176] <= 16'hFFFF;
rommem[12177] <= 16'hFFFF;
rommem[12178] <= 16'hFFFF;
rommem[12179] <= 16'hFFFF;
rommem[12180] <= 16'hFFFF;
rommem[12181] <= 16'hFFFF;
rommem[12182] <= 16'hFFFF;
rommem[12183] <= 16'hFFFF;
rommem[12184] <= 16'hFFFF;
rommem[12185] <= 16'hFFFF;
rommem[12186] <= 16'hFFFF;
rommem[12187] <= 16'hFFFF;
rommem[12188] <= 16'hFFFF;
rommem[12189] <= 16'hFFFF;
rommem[12190] <= 16'hFFFF;
rommem[12191] <= 16'hFFFF;
rommem[12192] <= 16'hFFFF;
rommem[12193] <= 16'hFFFF;
rommem[12194] <= 16'hFFFF;
rommem[12195] <= 16'hFFFF;
rommem[12196] <= 16'hFFFF;
rommem[12197] <= 16'hFFFF;
rommem[12198] <= 16'hFFFF;
rommem[12199] <= 16'hFFFF;
rommem[12200] <= 16'hFFFF;
rommem[12201] <= 16'hFFFF;
rommem[12202] <= 16'hFFFF;
rommem[12203] <= 16'hFFFF;
rommem[12204] <= 16'hFFFF;
rommem[12205] <= 16'hFFFF;
rommem[12206] <= 16'hFFFF;
rommem[12207] <= 16'hFFFF;
rommem[12208] <= 16'hFFFF;
rommem[12209] <= 16'hFFFF;
rommem[12210] <= 16'hFFFF;
rommem[12211] <= 16'hFFFF;
rommem[12212] <= 16'hFFFF;
rommem[12213] <= 16'hFFFF;
rommem[12214] <= 16'hFFFF;
rommem[12215] <= 16'hFFFF;
rommem[12216] <= 16'hFFFF;
rommem[12217] <= 16'hFFFF;
rommem[12218] <= 16'hFFFF;
rommem[12219] <= 16'hFFFF;
rommem[12220] <= 16'hFFFF;
rommem[12221] <= 16'hFFFF;
rommem[12222] <= 16'hFFFF;
rommem[12223] <= 16'hFFFF;
rommem[12224] <= 16'hFFFF;
rommem[12225] <= 16'hFFFF;
rommem[12226] <= 16'hFFFF;
rommem[12227] <= 16'hFFFF;
rommem[12228] <= 16'hFFFF;
rommem[12229] <= 16'hFFFF;
rommem[12230] <= 16'hFFFF;
rommem[12231] <= 16'hFFFF;
rommem[12232] <= 16'hFFFF;
rommem[12233] <= 16'hFFFF;
rommem[12234] <= 16'hFFFF;
rommem[12235] <= 16'hFFFF;
rommem[12236] <= 16'hFFFF;
rommem[12237] <= 16'hFFFF;
rommem[12238] <= 16'hFFFF;
rommem[12239] <= 16'hFFFF;
rommem[12240] <= 16'hFFFF;
rommem[12241] <= 16'hFFFF;
rommem[12242] <= 16'hFFFF;
rommem[12243] <= 16'hFFFF;
rommem[12244] <= 16'hFFFF;
rommem[12245] <= 16'hFFFF;
rommem[12246] <= 16'hFFFF;
rommem[12247] <= 16'hFFFF;
rommem[12248] <= 16'hFFFF;
rommem[12249] <= 16'hFFFF;
rommem[12250] <= 16'hFFFF;
rommem[12251] <= 16'hFFFF;
rommem[12252] <= 16'hFFFF;
rommem[12253] <= 16'hFFFF;
rommem[12254] <= 16'hFFFF;
rommem[12255] <= 16'hFFFF;
rommem[12256] <= 16'hFFFF;
rommem[12257] <= 16'hFFFF;
rommem[12258] <= 16'hFFFF;
rommem[12259] <= 16'hFFFF;
rommem[12260] <= 16'hFFFF;
rommem[12261] <= 16'hFFFF;
rommem[12262] <= 16'hFFFF;
rommem[12263] <= 16'hFFFF;
rommem[12264] <= 16'hFFFF;
rommem[12265] <= 16'hFFFF;
rommem[12266] <= 16'hFFFF;
rommem[12267] <= 16'hFFFF;
rommem[12268] <= 16'hFFFF;
rommem[12269] <= 16'hFFFF;
rommem[12270] <= 16'hFFFF;
rommem[12271] <= 16'hFFFF;
rommem[12272] <= 16'hFFFF;
rommem[12273] <= 16'hFFFF;
rommem[12274] <= 16'hFFFF;
rommem[12275] <= 16'hFFFF;
rommem[12276] <= 16'hFFFF;
rommem[12277] <= 16'hFFFF;
rommem[12278] <= 16'hFFFF;
rommem[12279] <= 16'hFFFF;
rommem[12280] <= 16'hFFFF;
rommem[12281] <= 16'hFFFF;
rommem[12282] <= 16'hFFFF;
rommem[12283] <= 16'hFFFF;
rommem[12284] <= 16'hFFFF;
rommem[12285] <= 16'hFFFF;
rommem[12286] <= 16'hFFFF;
rommem[12287] <= 16'hFFFF;
rommem[12288] <= 16'hFFFF;
rommem[12289] <= 16'hFFFF;
rommem[12290] <= 16'hFFFF;
rommem[12291] <= 16'hFFFF;
rommem[12292] <= 16'hFFFF;
rommem[12293] <= 16'hFFFF;
rommem[12294] <= 16'hFFFF;
rommem[12295] <= 16'hFFFF;
rommem[12296] <= 16'hFFFF;
rommem[12297] <= 16'hFFFF;
rommem[12298] <= 16'hFFFF;
rommem[12299] <= 16'hFFFF;
rommem[12300] <= 16'hFFFF;
rommem[12301] <= 16'hFFFF;
rommem[12302] <= 16'hFFFF;
rommem[12303] <= 16'hFFFF;
rommem[12304] <= 16'hFFFF;
rommem[12305] <= 16'hFFFF;
rommem[12306] <= 16'hFFFF;
rommem[12307] <= 16'hFFFF;
rommem[12308] <= 16'hFFFF;
rommem[12309] <= 16'hFFFF;
rommem[12310] <= 16'hFFFF;
rommem[12311] <= 16'hFFFF;
rommem[12312] <= 16'hFFFF;
rommem[12313] <= 16'hFFFF;
rommem[12314] <= 16'hFFFF;
rommem[12315] <= 16'hFFFF;
rommem[12316] <= 16'hFFFF;
rommem[12317] <= 16'hFFFF;
rommem[12318] <= 16'hFFFF;
rommem[12319] <= 16'hFFFF;
rommem[12320] <= 16'hFFFF;
rommem[12321] <= 16'hFFFF;
rommem[12322] <= 16'hFFFF;
rommem[12323] <= 16'hFFFF;
rommem[12324] <= 16'hFFFF;
rommem[12325] <= 16'hFFFF;
rommem[12326] <= 16'hFFFF;
rommem[12327] <= 16'hFFFF;
rommem[12328] <= 16'hFFFF;
rommem[12329] <= 16'hFFFF;
rommem[12330] <= 16'hFFFF;
rommem[12331] <= 16'hFFFF;
rommem[12332] <= 16'hFFFF;
rommem[12333] <= 16'hFFFF;
rommem[12334] <= 16'hFFFF;
rommem[12335] <= 16'hFFFF;
rommem[12336] <= 16'hFFFF;
rommem[12337] <= 16'hFFFF;
rommem[12338] <= 16'hFFFF;
rommem[12339] <= 16'hFFFF;
rommem[12340] <= 16'hFFFF;
rommem[12341] <= 16'hFFFF;
rommem[12342] <= 16'hFFFF;
rommem[12343] <= 16'hFFFF;
rommem[12344] <= 16'hFFFF;
rommem[12345] <= 16'hFFFF;
rommem[12346] <= 16'hFFFF;
rommem[12347] <= 16'hFFFF;
rommem[12348] <= 16'hFFFF;
rommem[12349] <= 16'hFFFF;
rommem[12350] <= 16'hFFFF;
rommem[12351] <= 16'hFFFF;
rommem[12352] <= 16'hFFFF;
rommem[12353] <= 16'hFFFF;
rommem[12354] <= 16'hFFFF;
rommem[12355] <= 16'hFFFF;
rommem[12356] <= 16'hFFFF;
rommem[12357] <= 16'hFFFF;
rommem[12358] <= 16'hFFFF;
rommem[12359] <= 16'hFFFF;
rommem[12360] <= 16'hFFFF;
rommem[12361] <= 16'hFFFF;
rommem[12362] <= 16'hFFFF;
rommem[12363] <= 16'hFFFF;
rommem[12364] <= 16'hFFFF;
rommem[12365] <= 16'hFFFF;
rommem[12366] <= 16'hFFFF;
rommem[12367] <= 16'hFFFF;
rommem[12368] <= 16'hFFFF;
rommem[12369] <= 16'hFFFF;
rommem[12370] <= 16'hFFFF;
rommem[12371] <= 16'hFFFF;
rommem[12372] <= 16'hFFFF;
rommem[12373] <= 16'hFFFF;
rommem[12374] <= 16'hFFFF;
rommem[12375] <= 16'hFFFF;
rommem[12376] <= 16'hFFFF;
rommem[12377] <= 16'hFFFF;
rommem[12378] <= 16'hFFFF;
rommem[12379] <= 16'hFFFF;
rommem[12380] <= 16'hFFFF;
rommem[12381] <= 16'hFFFF;
rommem[12382] <= 16'hFFFF;
rommem[12383] <= 16'hFFFF;
rommem[12384] <= 16'hFFFF;
rommem[12385] <= 16'hFFFF;
rommem[12386] <= 16'hFFFF;
rommem[12387] <= 16'hFFFF;
rommem[12388] <= 16'hFFFF;
rommem[12389] <= 16'hFFFF;
rommem[12390] <= 16'hFFFF;
rommem[12391] <= 16'hFFFF;
rommem[12392] <= 16'hFFFF;
rommem[12393] <= 16'hFFFF;
rommem[12394] <= 16'hFFFF;
rommem[12395] <= 16'hFFFF;
rommem[12396] <= 16'hFFFF;
rommem[12397] <= 16'hFFFF;
rommem[12398] <= 16'hFFFF;
rommem[12399] <= 16'hFFFF;
rommem[12400] <= 16'hFFFF;
rommem[12401] <= 16'hFFFF;
rommem[12402] <= 16'hFFFF;
rommem[12403] <= 16'hFFFF;
rommem[12404] <= 16'hFFFF;
rommem[12405] <= 16'hFFFF;
rommem[12406] <= 16'hFFFF;
rommem[12407] <= 16'hFFFF;
rommem[12408] <= 16'hFFFF;
rommem[12409] <= 16'hFFFF;
rommem[12410] <= 16'hFFFF;
rommem[12411] <= 16'hFFFF;
rommem[12412] <= 16'hFFFF;
rommem[12413] <= 16'hFFFF;
rommem[12414] <= 16'hFFFF;
rommem[12415] <= 16'hFFFF;
rommem[12416] <= 16'hFFFF;
rommem[12417] <= 16'hFFFF;
rommem[12418] <= 16'hFFFF;
rommem[12419] <= 16'hFFFF;
rommem[12420] <= 16'hFFFF;
rommem[12421] <= 16'hFFFF;
rommem[12422] <= 16'hFFFF;
rommem[12423] <= 16'hFFFF;
rommem[12424] <= 16'hFFFF;
rommem[12425] <= 16'hFFFF;
rommem[12426] <= 16'hFFFF;
rommem[12427] <= 16'hFFFF;
rommem[12428] <= 16'hFFFF;
rommem[12429] <= 16'hFFFF;
rommem[12430] <= 16'hFFFF;
rommem[12431] <= 16'hFFFF;
rommem[12432] <= 16'hFFFF;
rommem[12433] <= 16'hFFFF;
rommem[12434] <= 16'hFFFF;
rommem[12435] <= 16'hFFFF;
rommem[12436] <= 16'hFFFF;
rommem[12437] <= 16'hFFFF;
rommem[12438] <= 16'hFFFF;
rommem[12439] <= 16'hFFFF;
rommem[12440] <= 16'hFFFF;
rommem[12441] <= 16'hFFFF;
rommem[12442] <= 16'hFFFF;
rommem[12443] <= 16'hFFFF;
rommem[12444] <= 16'hFFFF;
rommem[12445] <= 16'hFFFF;
rommem[12446] <= 16'hFFFF;
rommem[12447] <= 16'hFFFF;
rommem[12448] <= 16'hFFFF;
rommem[12449] <= 16'hFFFF;
rommem[12450] <= 16'hFFFF;
rommem[12451] <= 16'hFFFF;
rommem[12452] <= 16'hFFFF;
rommem[12453] <= 16'hFFFF;
rommem[12454] <= 16'hFFFF;
rommem[12455] <= 16'hFFFF;
rommem[12456] <= 16'hFFFF;
rommem[12457] <= 16'hFFFF;
rommem[12458] <= 16'hFFFF;
rommem[12459] <= 16'hFFFF;
rommem[12460] <= 16'hFFFF;
rommem[12461] <= 16'hFFFF;
rommem[12462] <= 16'hFFFF;
rommem[12463] <= 16'hFFFF;
rommem[12464] <= 16'hFFFF;
rommem[12465] <= 16'hFFFF;
rommem[12466] <= 16'hFFFF;
rommem[12467] <= 16'hFFFF;
rommem[12468] <= 16'hFFFF;
rommem[12469] <= 16'hFFFF;
rommem[12470] <= 16'hFFFF;
rommem[12471] <= 16'hFFFF;
rommem[12472] <= 16'hFFFF;
rommem[12473] <= 16'hFFFF;
rommem[12474] <= 16'hFFFF;
rommem[12475] <= 16'hFFFF;
rommem[12476] <= 16'hFFFF;
rommem[12477] <= 16'hFFFF;
rommem[12478] <= 16'hFFFF;
rommem[12479] <= 16'hFFFF;
rommem[12480] <= 16'hFFFF;
rommem[12481] <= 16'hFFFF;
rommem[12482] <= 16'hFFFF;
rommem[12483] <= 16'hFFFF;
rommem[12484] <= 16'hFFFF;
rommem[12485] <= 16'hFFFF;
rommem[12486] <= 16'hFFFF;
rommem[12487] <= 16'hFFFF;
rommem[12488] <= 16'hFFFF;
rommem[12489] <= 16'hFFFF;
rommem[12490] <= 16'hFFFF;
rommem[12491] <= 16'hFFFF;
rommem[12492] <= 16'hFFFF;
rommem[12493] <= 16'hFFFF;
rommem[12494] <= 16'hFFFF;
rommem[12495] <= 16'hFFFF;
rommem[12496] <= 16'hFFFF;
rommem[12497] <= 16'hFFFF;
rommem[12498] <= 16'hFFFF;
rommem[12499] <= 16'hFFFF;
rommem[12500] <= 16'hFFFF;
rommem[12501] <= 16'hFFFF;
rommem[12502] <= 16'hFFFF;
rommem[12503] <= 16'hFFFF;
rommem[12504] <= 16'hFFFF;
rommem[12505] <= 16'hFFFF;
rommem[12506] <= 16'hFFFF;
rommem[12507] <= 16'hFFFF;
rommem[12508] <= 16'hFFFF;
rommem[12509] <= 16'hFFFF;
rommem[12510] <= 16'hFFFF;
rommem[12511] <= 16'hFFFF;
rommem[12512] <= 16'hFFFF;
rommem[12513] <= 16'hFFFF;
rommem[12514] <= 16'hFFFF;
rommem[12515] <= 16'hFFFF;
rommem[12516] <= 16'hFFFF;
rommem[12517] <= 16'hFFFF;
rommem[12518] <= 16'hFFFF;
rommem[12519] <= 16'hFFFF;
rommem[12520] <= 16'hFFFF;
rommem[12521] <= 16'hFFFF;
rommem[12522] <= 16'hFFFF;
rommem[12523] <= 16'hFFFF;
rommem[12524] <= 16'hFFFF;
rommem[12525] <= 16'hFFFF;
rommem[12526] <= 16'hFFFF;
rommem[12527] <= 16'hFFFF;
rommem[12528] <= 16'hFFFF;
rommem[12529] <= 16'hFFFF;
rommem[12530] <= 16'hFFFF;
rommem[12531] <= 16'hFFFF;
rommem[12532] <= 16'hFFFF;
rommem[12533] <= 16'hFFFF;
rommem[12534] <= 16'hFFFF;
rommem[12535] <= 16'hFFFF;
rommem[12536] <= 16'hFFFF;
rommem[12537] <= 16'hFFFF;
rommem[12538] <= 16'hFFFF;
rommem[12539] <= 16'hFFFF;
rommem[12540] <= 16'hFFFF;
rommem[12541] <= 16'hFFFF;
rommem[12542] <= 16'hFFFF;
rommem[12543] <= 16'hFFFF;
rommem[12544] <= 16'hFFFF;
rommem[12545] <= 16'hFFFF;
rommem[12546] <= 16'hFFFF;
rommem[12547] <= 16'hFFFF;
rommem[12548] <= 16'hFFFF;
rommem[12549] <= 16'hFFFF;
rommem[12550] <= 16'hFFFF;
rommem[12551] <= 16'hFFFF;
rommem[12552] <= 16'hFFFF;
rommem[12553] <= 16'hFFFF;
rommem[12554] <= 16'hFFFF;
rommem[12555] <= 16'hFFFF;
rommem[12556] <= 16'hFFFF;
rommem[12557] <= 16'hFFFF;
rommem[12558] <= 16'hFFFF;
rommem[12559] <= 16'hFFFF;
rommem[12560] <= 16'hFFFF;
rommem[12561] <= 16'hFFFF;
rommem[12562] <= 16'hFFFF;
rommem[12563] <= 16'hFFFF;
rommem[12564] <= 16'hFFFF;
rommem[12565] <= 16'hFFFF;
rommem[12566] <= 16'hFFFF;
rommem[12567] <= 16'hFFFF;
rommem[12568] <= 16'hFFFF;
rommem[12569] <= 16'hFFFF;
rommem[12570] <= 16'hFFFF;
rommem[12571] <= 16'hFFFF;
rommem[12572] <= 16'hFFFF;
rommem[12573] <= 16'hFFFF;
rommem[12574] <= 16'hFFFF;
rommem[12575] <= 16'hFFFF;
rommem[12576] <= 16'hFFFF;
rommem[12577] <= 16'hFFFF;
rommem[12578] <= 16'hFFFF;
rommem[12579] <= 16'hFFFF;
rommem[12580] <= 16'hFFFF;
rommem[12581] <= 16'hFFFF;
rommem[12582] <= 16'hFFFF;
rommem[12583] <= 16'hFFFF;
rommem[12584] <= 16'hFFFF;
rommem[12585] <= 16'hFFFF;
rommem[12586] <= 16'hFFFF;
rommem[12587] <= 16'hFFFF;
rommem[12588] <= 16'hFFFF;
rommem[12589] <= 16'hFFFF;
rommem[12590] <= 16'hFFFF;
rommem[12591] <= 16'hFFFF;
rommem[12592] <= 16'hFFFF;
rommem[12593] <= 16'hFFFF;
rommem[12594] <= 16'hFFFF;
rommem[12595] <= 16'hFFFF;
rommem[12596] <= 16'hFFFF;
rommem[12597] <= 16'hFFFF;
rommem[12598] <= 16'hFFFF;
rommem[12599] <= 16'hFFFF;
rommem[12600] <= 16'hFFFF;
rommem[12601] <= 16'hFFFF;
rommem[12602] <= 16'hFFFF;
rommem[12603] <= 16'hFFFF;
rommem[12604] <= 16'hFFFF;
rommem[12605] <= 16'hFFFF;
rommem[12606] <= 16'hFFFF;
rommem[12607] <= 16'hFFFF;
rommem[12608] <= 16'hFFFF;
rommem[12609] <= 16'hFFFF;
rommem[12610] <= 16'hFFFF;
rommem[12611] <= 16'hFFFF;
rommem[12612] <= 16'hFFFF;
rommem[12613] <= 16'hFFFF;
rommem[12614] <= 16'hFFFF;
rommem[12615] <= 16'hFFFF;
rommem[12616] <= 16'hFFFF;
rommem[12617] <= 16'hFFFF;
rommem[12618] <= 16'hFFFF;
rommem[12619] <= 16'hFFFF;
rommem[12620] <= 16'hFFFF;
rommem[12621] <= 16'hFFFF;
rommem[12622] <= 16'hFFFF;
rommem[12623] <= 16'hFFFF;
rommem[12624] <= 16'hFFFF;
rommem[12625] <= 16'hFFFF;
rommem[12626] <= 16'hFFFF;
rommem[12627] <= 16'hFFFF;
rommem[12628] <= 16'hFFFF;
rommem[12629] <= 16'hFFFF;
rommem[12630] <= 16'hFFFF;
rommem[12631] <= 16'hFFFF;
rommem[12632] <= 16'hFFFF;
rommem[12633] <= 16'hFFFF;
rommem[12634] <= 16'hFFFF;
rommem[12635] <= 16'hFFFF;
rommem[12636] <= 16'hFFFF;
rommem[12637] <= 16'hFFFF;
rommem[12638] <= 16'hFFFF;
rommem[12639] <= 16'hFFFF;
rommem[12640] <= 16'hFFFF;
rommem[12641] <= 16'hFFFF;
rommem[12642] <= 16'hFFFF;
rommem[12643] <= 16'hFFFF;
rommem[12644] <= 16'hFFFF;
rommem[12645] <= 16'hFFFF;
rommem[12646] <= 16'hFFFF;
rommem[12647] <= 16'hFFFF;
rommem[12648] <= 16'hFFFF;
rommem[12649] <= 16'hFFFF;
rommem[12650] <= 16'hFFFF;
rommem[12651] <= 16'hFFFF;
rommem[12652] <= 16'hFFFF;
rommem[12653] <= 16'hFFFF;
rommem[12654] <= 16'hFFFF;
rommem[12655] <= 16'hFFFF;
rommem[12656] <= 16'hFFFF;
rommem[12657] <= 16'hFFFF;
rommem[12658] <= 16'hFFFF;
rommem[12659] <= 16'hFFFF;
rommem[12660] <= 16'hFFFF;
rommem[12661] <= 16'hFFFF;
rommem[12662] <= 16'hFFFF;
rommem[12663] <= 16'hFFFF;
rommem[12664] <= 16'hFFFF;
rommem[12665] <= 16'hFFFF;
rommem[12666] <= 16'hFFFF;
rommem[12667] <= 16'hFFFF;
rommem[12668] <= 16'hFFFF;
rommem[12669] <= 16'hFFFF;
rommem[12670] <= 16'hFFFF;
rommem[12671] <= 16'hFFFF;
rommem[12672] <= 16'hFFFF;
rommem[12673] <= 16'hFFFF;
rommem[12674] <= 16'hFFFF;
rommem[12675] <= 16'hFFFF;
rommem[12676] <= 16'hFFFF;
rommem[12677] <= 16'hFFFF;
rommem[12678] <= 16'hFFFF;
rommem[12679] <= 16'hFFFF;
rommem[12680] <= 16'hFFFF;
rommem[12681] <= 16'hFFFF;
rommem[12682] <= 16'hFFFF;
rommem[12683] <= 16'hFFFF;
rommem[12684] <= 16'hFFFF;
rommem[12685] <= 16'hFFFF;
rommem[12686] <= 16'hFFFF;
rommem[12687] <= 16'hFFFF;
rommem[12688] <= 16'hFFFF;
rommem[12689] <= 16'hFFFF;
rommem[12690] <= 16'hFFFF;
rommem[12691] <= 16'hFFFF;
rommem[12692] <= 16'hFFFF;
rommem[12693] <= 16'hFFFF;
rommem[12694] <= 16'hFFFF;
rommem[12695] <= 16'hFFFF;
rommem[12696] <= 16'hFFFF;
rommem[12697] <= 16'hFFFF;
rommem[12698] <= 16'hFFFF;
rommem[12699] <= 16'hFFFF;
rommem[12700] <= 16'hFFFF;
rommem[12701] <= 16'hFFFF;
rommem[12702] <= 16'hFFFF;
rommem[12703] <= 16'hFFFF;
rommem[12704] <= 16'hFFFF;
rommem[12705] <= 16'hFFFF;
rommem[12706] <= 16'hFFFF;
rommem[12707] <= 16'hFFFF;
rommem[12708] <= 16'hFFFF;
rommem[12709] <= 16'hFFFF;
rommem[12710] <= 16'hFFFF;
rommem[12711] <= 16'hFFFF;
rommem[12712] <= 16'hFFFF;
rommem[12713] <= 16'hFFFF;
rommem[12714] <= 16'hFFFF;
rommem[12715] <= 16'hFFFF;
rommem[12716] <= 16'hFFFF;
rommem[12717] <= 16'hFFFF;
rommem[12718] <= 16'hFFFF;
rommem[12719] <= 16'hFFFF;
rommem[12720] <= 16'hFFFF;
rommem[12721] <= 16'hFFFF;
rommem[12722] <= 16'hFFFF;
rommem[12723] <= 16'hFFFF;
rommem[12724] <= 16'hFFFF;
rommem[12725] <= 16'hFFFF;
rommem[12726] <= 16'hFFFF;
rommem[12727] <= 16'hFFFF;
rommem[12728] <= 16'hFFFF;
rommem[12729] <= 16'hFFFF;
rommem[12730] <= 16'hFFFF;
rommem[12731] <= 16'hFFFF;
rommem[12732] <= 16'hFFFF;
rommem[12733] <= 16'hFFFF;
rommem[12734] <= 16'hFFFF;
rommem[12735] <= 16'hFFFF;
rommem[12736] <= 16'hFFFF;
rommem[12737] <= 16'hFFFF;
rommem[12738] <= 16'hFFFF;
rommem[12739] <= 16'hFFFF;
rommem[12740] <= 16'hFFFF;
rommem[12741] <= 16'hFFFF;
rommem[12742] <= 16'hFFFF;
rommem[12743] <= 16'hFFFF;
rommem[12744] <= 16'hFFFF;
rommem[12745] <= 16'hFFFF;
rommem[12746] <= 16'hFFFF;
rommem[12747] <= 16'hFFFF;
rommem[12748] <= 16'hFFFF;
rommem[12749] <= 16'hFFFF;
rommem[12750] <= 16'hFFFF;
rommem[12751] <= 16'hFFFF;
rommem[12752] <= 16'hFFFF;
rommem[12753] <= 16'hFFFF;
rommem[12754] <= 16'hFFFF;
rommem[12755] <= 16'hFFFF;
rommem[12756] <= 16'hFFFF;
rommem[12757] <= 16'hFFFF;
rommem[12758] <= 16'hFFFF;
rommem[12759] <= 16'hFFFF;
rommem[12760] <= 16'hFFFF;
rommem[12761] <= 16'hFFFF;
rommem[12762] <= 16'hFFFF;
rommem[12763] <= 16'hFFFF;
rommem[12764] <= 16'hFFFF;
rommem[12765] <= 16'hFFFF;
rommem[12766] <= 16'hFFFF;
rommem[12767] <= 16'hFFFF;
rommem[12768] <= 16'hFFFF;
rommem[12769] <= 16'hFFFF;
rommem[12770] <= 16'hFFFF;
rommem[12771] <= 16'hFFFF;
rommem[12772] <= 16'hFFFF;
rommem[12773] <= 16'hFFFF;
rommem[12774] <= 16'hFFFF;
rommem[12775] <= 16'hFFFF;
rommem[12776] <= 16'hFFFF;
rommem[12777] <= 16'hFFFF;
rommem[12778] <= 16'hFFFF;
rommem[12779] <= 16'hFFFF;
rommem[12780] <= 16'hFFFF;
rommem[12781] <= 16'hFFFF;
rommem[12782] <= 16'hFFFF;
rommem[12783] <= 16'hFFFF;
rommem[12784] <= 16'hFFFF;
rommem[12785] <= 16'hFFFF;
rommem[12786] <= 16'hFFFF;
rommem[12787] <= 16'hFFFF;
rommem[12788] <= 16'hFFFF;
rommem[12789] <= 16'hFFFF;
rommem[12790] <= 16'hFFFF;
rommem[12791] <= 16'hFFFF;
rommem[12792] <= 16'hFFFF;
rommem[12793] <= 16'hFFFF;
rommem[12794] <= 16'hFFFF;
rommem[12795] <= 16'hFFFF;
rommem[12796] <= 16'hFFFF;
rommem[12797] <= 16'hFFFF;
rommem[12798] <= 16'hFFFF;
rommem[12799] <= 16'hFFFF;
rommem[12800] <= 16'hFFFF;
rommem[12801] <= 16'hFFFF;
rommem[12802] <= 16'hFFFF;
rommem[12803] <= 16'hFFFF;
rommem[12804] <= 16'hFFFF;
rommem[12805] <= 16'hFFFF;
rommem[12806] <= 16'hFFFF;
rommem[12807] <= 16'hFFFF;
rommem[12808] <= 16'hFFFF;
rommem[12809] <= 16'hFFFF;
rommem[12810] <= 16'hFFFF;
rommem[12811] <= 16'hFFFF;
rommem[12812] <= 16'hFFFF;
rommem[12813] <= 16'hFFFF;
rommem[12814] <= 16'hFFFF;
rommem[12815] <= 16'hFFFF;
rommem[12816] <= 16'hFFFF;
rommem[12817] <= 16'hFFFF;
rommem[12818] <= 16'hFFFF;
rommem[12819] <= 16'hFFFF;
rommem[12820] <= 16'hFFFF;
rommem[12821] <= 16'hFFFF;
rommem[12822] <= 16'hFFFF;
rommem[12823] <= 16'hFFFF;
rommem[12824] <= 16'hFFFF;
rommem[12825] <= 16'hFFFF;
rommem[12826] <= 16'hFFFF;
rommem[12827] <= 16'hFFFF;
rommem[12828] <= 16'hFFFF;
rommem[12829] <= 16'hFFFF;
rommem[12830] <= 16'hFFFF;
rommem[12831] <= 16'hFFFF;
rommem[12832] <= 16'hFFFF;
rommem[12833] <= 16'hFFFF;
rommem[12834] <= 16'hFFFF;
rommem[12835] <= 16'hFFFF;
rommem[12836] <= 16'hFFFF;
rommem[12837] <= 16'hFFFF;
rommem[12838] <= 16'hFFFF;
rommem[12839] <= 16'hFFFF;
rommem[12840] <= 16'hFFFF;
rommem[12841] <= 16'hFFFF;
rommem[12842] <= 16'hFFFF;
rommem[12843] <= 16'hFFFF;
rommem[12844] <= 16'hFFFF;
rommem[12845] <= 16'hFFFF;
rommem[12846] <= 16'hFFFF;
rommem[12847] <= 16'hFFFF;
rommem[12848] <= 16'hFFFF;
rommem[12849] <= 16'hFFFF;
rommem[12850] <= 16'hFFFF;
rommem[12851] <= 16'hFFFF;
rommem[12852] <= 16'hFFFF;
rommem[12853] <= 16'hFFFF;
rommem[12854] <= 16'hFFFF;
rommem[12855] <= 16'hFFFF;
rommem[12856] <= 16'hFFFF;
rommem[12857] <= 16'hFFFF;
rommem[12858] <= 16'hFFFF;
rommem[12859] <= 16'hFFFF;
rommem[12860] <= 16'hFFFF;
rommem[12861] <= 16'hFFFF;
rommem[12862] <= 16'hFFFF;
rommem[12863] <= 16'hFFFF;
rommem[12864] <= 16'hFFFF;
rommem[12865] <= 16'hFFFF;
rommem[12866] <= 16'hFFFF;
rommem[12867] <= 16'hFFFF;
rommem[12868] <= 16'hFFFF;
rommem[12869] <= 16'hFFFF;
rommem[12870] <= 16'hFFFF;
rommem[12871] <= 16'hFFFF;
rommem[12872] <= 16'hFFFF;
rommem[12873] <= 16'hFFFF;
rommem[12874] <= 16'hFFFF;
rommem[12875] <= 16'hFFFF;
rommem[12876] <= 16'hFFFF;
rommem[12877] <= 16'hFFFF;
rommem[12878] <= 16'hFFFF;
rommem[12879] <= 16'hFFFF;
rommem[12880] <= 16'hFFFF;
rommem[12881] <= 16'hFFFF;
rommem[12882] <= 16'hFFFF;
rommem[12883] <= 16'hFFFF;
rommem[12884] <= 16'hFFFF;
rommem[12885] <= 16'hFFFF;
rommem[12886] <= 16'hFFFF;
rommem[12887] <= 16'hFFFF;
rommem[12888] <= 16'hFFFF;
rommem[12889] <= 16'hFFFF;
rommem[12890] <= 16'hFFFF;
rommem[12891] <= 16'hFFFF;
rommem[12892] <= 16'hFFFF;
rommem[12893] <= 16'hFFFF;
rommem[12894] <= 16'hFFFF;
rommem[12895] <= 16'hFFFF;
rommem[12896] <= 16'hFFFF;
rommem[12897] <= 16'hFFFF;
rommem[12898] <= 16'hFFFF;
rommem[12899] <= 16'hFFFF;
rommem[12900] <= 16'hFFFF;
rommem[12901] <= 16'hFFFF;
rommem[12902] <= 16'hFFFF;
rommem[12903] <= 16'hFFFF;
rommem[12904] <= 16'hFFFF;
rommem[12905] <= 16'hFFFF;
rommem[12906] <= 16'hFFFF;
rommem[12907] <= 16'hFFFF;
rommem[12908] <= 16'hFFFF;
rommem[12909] <= 16'hFFFF;
rommem[12910] <= 16'hFFFF;
rommem[12911] <= 16'hFFFF;
rommem[12912] <= 16'hFFFF;
rommem[12913] <= 16'hFFFF;
rommem[12914] <= 16'hFFFF;
rommem[12915] <= 16'hFFFF;
rommem[12916] <= 16'hFFFF;
rommem[12917] <= 16'hFFFF;
rommem[12918] <= 16'hFFFF;
rommem[12919] <= 16'hFFFF;
rommem[12920] <= 16'hFFFF;
rommem[12921] <= 16'hFFFF;
rommem[12922] <= 16'hFFFF;
rommem[12923] <= 16'hFFFF;
rommem[12924] <= 16'hFFFF;
rommem[12925] <= 16'hFFFF;
rommem[12926] <= 16'hFFFF;
rommem[12927] <= 16'hFFFF;
rommem[12928] <= 16'hFFFF;
rommem[12929] <= 16'hFFFF;
rommem[12930] <= 16'hFFFF;
rommem[12931] <= 16'hFFFF;
rommem[12932] <= 16'hFFFF;
rommem[12933] <= 16'hFFFF;
rommem[12934] <= 16'hFFFF;
rommem[12935] <= 16'hFFFF;
rommem[12936] <= 16'hFFFF;
rommem[12937] <= 16'hFFFF;
rommem[12938] <= 16'hFFFF;
rommem[12939] <= 16'hFFFF;
rommem[12940] <= 16'hFFFF;
rommem[12941] <= 16'hFFFF;
rommem[12942] <= 16'hFFFF;
rommem[12943] <= 16'hFFFF;
rommem[12944] <= 16'hFFFF;
rommem[12945] <= 16'hFFFF;
rommem[12946] <= 16'hFFFF;
rommem[12947] <= 16'hFFFF;
rommem[12948] <= 16'hFFFF;
rommem[12949] <= 16'hFFFF;
rommem[12950] <= 16'hFFFF;
rommem[12951] <= 16'hFFFF;
rommem[12952] <= 16'hFFFF;
rommem[12953] <= 16'hFFFF;
rommem[12954] <= 16'hFFFF;
rommem[12955] <= 16'hFFFF;
rommem[12956] <= 16'hFFFF;
rommem[12957] <= 16'hFFFF;
rommem[12958] <= 16'hFFFF;
rommem[12959] <= 16'hFFFF;
rommem[12960] <= 16'hFFFF;
rommem[12961] <= 16'hFFFF;
rommem[12962] <= 16'hFFFF;
rommem[12963] <= 16'hFFFF;
rommem[12964] <= 16'hFFFF;
rommem[12965] <= 16'hFFFF;
rommem[12966] <= 16'hFFFF;
rommem[12967] <= 16'hFFFF;
rommem[12968] <= 16'hFFFF;
rommem[12969] <= 16'hFFFF;
rommem[12970] <= 16'hFFFF;
rommem[12971] <= 16'hFFFF;
rommem[12972] <= 16'hFFFF;
rommem[12973] <= 16'hFFFF;
rommem[12974] <= 16'hFFFF;
rommem[12975] <= 16'hFFFF;
rommem[12976] <= 16'hFFFF;
rommem[12977] <= 16'hFFFF;
rommem[12978] <= 16'hFFFF;
rommem[12979] <= 16'hFFFF;
rommem[12980] <= 16'hFFFF;
rommem[12981] <= 16'hFFFF;
rommem[12982] <= 16'hFFFF;
rommem[12983] <= 16'hFFFF;
rommem[12984] <= 16'hFFFF;
rommem[12985] <= 16'hFFFF;
rommem[12986] <= 16'hFFFF;
rommem[12987] <= 16'hFFFF;
rommem[12988] <= 16'hFFFF;
rommem[12989] <= 16'hFFFF;
rommem[12990] <= 16'hFFFF;
rommem[12991] <= 16'hFFFF;
rommem[12992] <= 16'hFFFF;
rommem[12993] <= 16'hFFFF;
rommem[12994] <= 16'hFFFF;
rommem[12995] <= 16'hFFFF;
rommem[12996] <= 16'hFFFF;
rommem[12997] <= 16'hFFFF;
rommem[12998] <= 16'hFFFF;
rommem[12999] <= 16'hFFFF;
rommem[13000] <= 16'hFFFF;
rommem[13001] <= 16'hFFFF;
rommem[13002] <= 16'hFFFF;
rommem[13003] <= 16'hFFFF;
rommem[13004] <= 16'hFFFF;
rommem[13005] <= 16'hFFFF;
rommem[13006] <= 16'hFFFF;
rommem[13007] <= 16'hFFFF;
rommem[13008] <= 16'hFFFF;
rommem[13009] <= 16'hFFFF;
rommem[13010] <= 16'hFFFF;
rommem[13011] <= 16'hFFFF;
rommem[13012] <= 16'hFFFF;
rommem[13013] <= 16'hFFFF;
rommem[13014] <= 16'hFFFF;
rommem[13015] <= 16'hFFFF;
rommem[13016] <= 16'hFFFF;
rommem[13017] <= 16'hFFFF;
rommem[13018] <= 16'hFFFF;
rommem[13019] <= 16'hFFFF;
rommem[13020] <= 16'hFFFF;
rommem[13021] <= 16'hFFFF;
rommem[13022] <= 16'hFFFF;
rommem[13023] <= 16'hFFFF;
rommem[13024] <= 16'hFFFF;
rommem[13025] <= 16'hFFFF;
rommem[13026] <= 16'hFFFF;
rommem[13027] <= 16'hFFFF;
rommem[13028] <= 16'hFFFF;
rommem[13029] <= 16'hFFFF;
rommem[13030] <= 16'hFFFF;
rommem[13031] <= 16'hFFFF;
rommem[13032] <= 16'hFFFF;
rommem[13033] <= 16'hFFFF;
rommem[13034] <= 16'hFFFF;
rommem[13035] <= 16'hFFFF;
rommem[13036] <= 16'hFFFF;
rommem[13037] <= 16'hFFFF;
rommem[13038] <= 16'hFFFF;
rommem[13039] <= 16'hFFFF;
rommem[13040] <= 16'hFFFF;
rommem[13041] <= 16'hFFFF;
rommem[13042] <= 16'hFFFF;
rommem[13043] <= 16'hFFFF;
rommem[13044] <= 16'hFFFF;
rommem[13045] <= 16'hFFFF;
rommem[13046] <= 16'hFFFF;
rommem[13047] <= 16'hFFFF;
rommem[13048] <= 16'hFFFF;
rommem[13049] <= 16'hFFFF;
rommem[13050] <= 16'hFFFF;
rommem[13051] <= 16'hFFFF;
rommem[13052] <= 16'hFFFF;
rommem[13053] <= 16'hFFFF;
rommem[13054] <= 16'hFFFF;
rommem[13055] <= 16'hFFFF;
rommem[13056] <= 16'hFFFF;
rommem[13057] <= 16'hFFFF;
rommem[13058] <= 16'hFFFF;
rommem[13059] <= 16'hFFFF;
rommem[13060] <= 16'hFFFF;
rommem[13061] <= 16'hFFFF;
rommem[13062] <= 16'hFFFF;
rommem[13063] <= 16'hFFFF;
rommem[13064] <= 16'hFFFF;
rommem[13065] <= 16'hFFFF;
rommem[13066] <= 16'hFFFF;
rommem[13067] <= 16'hFFFF;
rommem[13068] <= 16'hFFFF;
rommem[13069] <= 16'hFFFF;
rommem[13070] <= 16'hFFFF;
rommem[13071] <= 16'hFFFF;
rommem[13072] <= 16'hFFFF;
rommem[13073] <= 16'hFFFF;
rommem[13074] <= 16'hFFFF;
rommem[13075] <= 16'hFFFF;
rommem[13076] <= 16'hFFFF;
rommem[13077] <= 16'hFFFF;
rommem[13078] <= 16'hFFFF;
rommem[13079] <= 16'hFFFF;
rommem[13080] <= 16'hFFFF;
rommem[13081] <= 16'hFFFF;
rommem[13082] <= 16'hFFFF;
rommem[13083] <= 16'hFFFF;
rommem[13084] <= 16'hFFFF;
rommem[13085] <= 16'hFFFF;
rommem[13086] <= 16'hFFFF;
rommem[13087] <= 16'hFFFF;
rommem[13088] <= 16'hFFFF;
rommem[13089] <= 16'hFFFF;
rommem[13090] <= 16'hFFFF;
rommem[13091] <= 16'hFFFF;
rommem[13092] <= 16'hFFFF;
rommem[13093] <= 16'hFFFF;
rommem[13094] <= 16'hFFFF;
rommem[13095] <= 16'hFFFF;
rommem[13096] <= 16'hFFFF;
rommem[13097] <= 16'hFFFF;
rommem[13098] <= 16'hFFFF;
rommem[13099] <= 16'hFFFF;
rommem[13100] <= 16'hFFFF;
rommem[13101] <= 16'hFFFF;
rommem[13102] <= 16'hFFFF;
rommem[13103] <= 16'hFFFF;
rommem[13104] <= 16'hFFFF;
rommem[13105] <= 16'hFFFF;
rommem[13106] <= 16'hFFFF;
rommem[13107] <= 16'hFFFF;
rommem[13108] <= 16'hFFFF;
rommem[13109] <= 16'hFFFF;
rommem[13110] <= 16'hFFFF;
rommem[13111] <= 16'hFFFF;
rommem[13112] <= 16'hFFFF;
rommem[13113] <= 16'hFFFF;
rommem[13114] <= 16'hFFFF;
rommem[13115] <= 16'hFFFF;
rommem[13116] <= 16'hFFFF;
rommem[13117] <= 16'hFFFF;
rommem[13118] <= 16'hFFFF;
rommem[13119] <= 16'hFFFF;
rommem[13120] <= 16'hFFFF;
rommem[13121] <= 16'hFFFF;
rommem[13122] <= 16'hFFFF;
rommem[13123] <= 16'hFFFF;
rommem[13124] <= 16'hFFFF;
rommem[13125] <= 16'hFFFF;
rommem[13126] <= 16'hFFFF;
rommem[13127] <= 16'hFFFF;
rommem[13128] <= 16'hFFFF;
rommem[13129] <= 16'hFFFF;
rommem[13130] <= 16'hFFFF;
rommem[13131] <= 16'hFFFF;
rommem[13132] <= 16'hFFFF;
rommem[13133] <= 16'hFFFF;
rommem[13134] <= 16'hFFFF;
rommem[13135] <= 16'hFFFF;
rommem[13136] <= 16'hFFFF;
rommem[13137] <= 16'hFFFF;
rommem[13138] <= 16'hFFFF;
rommem[13139] <= 16'hFFFF;
rommem[13140] <= 16'hFFFF;
rommem[13141] <= 16'hFFFF;
rommem[13142] <= 16'hFFFF;
rommem[13143] <= 16'hFFFF;
rommem[13144] <= 16'hFFFF;
rommem[13145] <= 16'hFFFF;
rommem[13146] <= 16'hFFFF;
rommem[13147] <= 16'hFFFF;
rommem[13148] <= 16'hFFFF;
rommem[13149] <= 16'hFFFF;
rommem[13150] <= 16'hFFFF;
rommem[13151] <= 16'hFFFF;
rommem[13152] <= 16'hFFFF;
rommem[13153] <= 16'hFFFF;
rommem[13154] <= 16'hFFFF;
rommem[13155] <= 16'hFFFF;
rommem[13156] <= 16'hFFFF;
rommem[13157] <= 16'hFFFF;
rommem[13158] <= 16'hFFFF;
rommem[13159] <= 16'hFFFF;
rommem[13160] <= 16'hFFFF;
rommem[13161] <= 16'hFFFF;
rommem[13162] <= 16'hFFFF;
rommem[13163] <= 16'hFFFF;
rommem[13164] <= 16'hFFFF;
rommem[13165] <= 16'hFFFF;
rommem[13166] <= 16'hFFFF;
rommem[13167] <= 16'hFFFF;
rommem[13168] <= 16'hFFFF;
rommem[13169] <= 16'hFFFF;
rommem[13170] <= 16'hFFFF;
rommem[13171] <= 16'hFFFF;
rommem[13172] <= 16'hFFFF;
rommem[13173] <= 16'hFFFF;
rommem[13174] <= 16'hFFFF;
rommem[13175] <= 16'hFFFF;
rommem[13176] <= 16'hFFFF;
rommem[13177] <= 16'hFFFF;
rommem[13178] <= 16'hFFFF;
rommem[13179] <= 16'hFFFF;
rommem[13180] <= 16'hFFFF;
rommem[13181] <= 16'hFFFF;
rommem[13182] <= 16'hFFFF;
rommem[13183] <= 16'hFFFF;
rommem[13184] <= 16'hFFFF;
rommem[13185] <= 16'hFFFF;
rommem[13186] <= 16'hFFFF;
rommem[13187] <= 16'hFFFF;
rommem[13188] <= 16'hFFFF;
rommem[13189] <= 16'hFFFF;
rommem[13190] <= 16'hFFFF;
rommem[13191] <= 16'hFFFF;
rommem[13192] <= 16'hFFFF;
rommem[13193] <= 16'hFFFF;
rommem[13194] <= 16'hFFFF;
rommem[13195] <= 16'hFFFF;
rommem[13196] <= 16'hFFFF;
rommem[13197] <= 16'hFFFF;
rommem[13198] <= 16'hFFFF;
rommem[13199] <= 16'hFFFF;
rommem[13200] <= 16'hFFFF;
rommem[13201] <= 16'hFFFF;
rommem[13202] <= 16'hFFFF;
rommem[13203] <= 16'hFFFF;
rommem[13204] <= 16'hFFFF;
rommem[13205] <= 16'hFFFF;
rommem[13206] <= 16'hFFFF;
rommem[13207] <= 16'hFFFF;
rommem[13208] <= 16'hFFFF;
rommem[13209] <= 16'hFFFF;
rommem[13210] <= 16'hFFFF;
rommem[13211] <= 16'hFFFF;
rommem[13212] <= 16'hFFFF;
rommem[13213] <= 16'hFFFF;
rommem[13214] <= 16'hFFFF;
rommem[13215] <= 16'hFFFF;
rommem[13216] <= 16'hFFFF;
rommem[13217] <= 16'hFFFF;
rommem[13218] <= 16'hFFFF;
rommem[13219] <= 16'hFFFF;
rommem[13220] <= 16'hFFFF;
rommem[13221] <= 16'hFFFF;
rommem[13222] <= 16'hFFFF;
rommem[13223] <= 16'hFFFF;
rommem[13224] <= 16'hFFFF;
rommem[13225] <= 16'hFFFF;
rommem[13226] <= 16'hFFFF;
rommem[13227] <= 16'hFFFF;
rommem[13228] <= 16'hFFFF;
rommem[13229] <= 16'hFFFF;
rommem[13230] <= 16'hFFFF;
rommem[13231] <= 16'hFFFF;
rommem[13232] <= 16'hFFFF;
rommem[13233] <= 16'hFFFF;
rommem[13234] <= 16'hFFFF;
rommem[13235] <= 16'hFFFF;
rommem[13236] <= 16'hFFFF;
rommem[13237] <= 16'hFFFF;
rommem[13238] <= 16'hFFFF;
rommem[13239] <= 16'hFFFF;
rommem[13240] <= 16'hFFFF;
rommem[13241] <= 16'hFFFF;
rommem[13242] <= 16'hFFFF;
rommem[13243] <= 16'hFFFF;
rommem[13244] <= 16'hFFFF;
rommem[13245] <= 16'hFFFF;
rommem[13246] <= 16'hFFFF;
rommem[13247] <= 16'hFFFF;
rommem[13248] <= 16'hFFFF;
rommem[13249] <= 16'hFFFF;
rommem[13250] <= 16'hFFFF;
rommem[13251] <= 16'hFFFF;
rommem[13252] <= 16'hFFFF;
rommem[13253] <= 16'hFFFF;
rommem[13254] <= 16'hFFFF;
rommem[13255] <= 16'hFFFF;
rommem[13256] <= 16'hFFFF;
rommem[13257] <= 16'hFFFF;
rommem[13258] <= 16'hFFFF;
rommem[13259] <= 16'hFFFF;
rommem[13260] <= 16'hFFFF;
rommem[13261] <= 16'hFFFF;
rommem[13262] <= 16'hFFFF;
rommem[13263] <= 16'hFFFF;
rommem[13264] <= 16'hFFFF;
rommem[13265] <= 16'hFFFF;
rommem[13266] <= 16'hFFFF;
rommem[13267] <= 16'hFFFF;
rommem[13268] <= 16'hFFFF;
rommem[13269] <= 16'hFFFF;
rommem[13270] <= 16'hFFFF;
rommem[13271] <= 16'hFFFF;
rommem[13272] <= 16'hFFFF;
rommem[13273] <= 16'hFFFF;
rommem[13274] <= 16'hFFFF;
rommem[13275] <= 16'hFFFF;
rommem[13276] <= 16'hFFFF;
rommem[13277] <= 16'hFFFF;
rommem[13278] <= 16'hFFFF;
rommem[13279] <= 16'hFFFF;
rommem[13280] <= 16'hFFFF;
rommem[13281] <= 16'hFFFF;
rommem[13282] <= 16'hFFFF;
rommem[13283] <= 16'hFFFF;
rommem[13284] <= 16'hFFFF;
rommem[13285] <= 16'hFFFF;
rommem[13286] <= 16'hFFFF;
rommem[13287] <= 16'hFFFF;
rommem[13288] <= 16'hFFFF;
rommem[13289] <= 16'hFFFF;
rommem[13290] <= 16'hFFFF;
rommem[13291] <= 16'hFFFF;
rommem[13292] <= 16'hFFFF;
rommem[13293] <= 16'hFFFF;
rommem[13294] <= 16'hFFFF;
rommem[13295] <= 16'hFFFF;
rommem[13296] <= 16'hFFFF;
rommem[13297] <= 16'hFFFF;
rommem[13298] <= 16'hFFFF;
rommem[13299] <= 16'hFFFF;
rommem[13300] <= 16'hFFFF;
rommem[13301] <= 16'hFFFF;
rommem[13302] <= 16'hFFFF;
rommem[13303] <= 16'hFFFF;
rommem[13304] <= 16'hFFFF;
rommem[13305] <= 16'hFFFF;
rommem[13306] <= 16'hFFFF;
rommem[13307] <= 16'hFFFF;
rommem[13308] <= 16'hFFFF;
rommem[13309] <= 16'hFFFF;
rommem[13310] <= 16'hFFFF;
rommem[13311] <= 16'hFFFF;
rommem[13312] <= 16'hFFFF;
rommem[13313] <= 16'hFFFF;
rommem[13314] <= 16'hFFFF;
rommem[13315] <= 16'hFFFF;
rommem[13316] <= 16'hFFFF;
rommem[13317] <= 16'hFFFF;
rommem[13318] <= 16'hFFFF;
rommem[13319] <= 16'hFFFF;
rommem[13320] <= 16'hFFFF;
rommem[13321] <= 16'hFFFF;
rommem[13322] <= 16'hFFFF;
rommem[13323] <= 16'hFFFF;
rommem[13324] <= 16'hFFFF;
rommem[13325] <= 16'hFFFF;
rommem[13326] <= 16'hFFFF;
rommem[13327] <= 16'hFFFF;
rommem[13328] <= 16'hFFFF;
rommem[13329] <= 16'hFFFF;
rommem[13330] <= 16'hFFFF;
rommem[13331] <= 16'hFFFF;
rommem[13332] <= 16'hFFFF;
rommem[13333] <= 16'hFFFF;
rommem[13334] <= 16'hFFFF;
rommem[13335] <= 16'hFFFF;
rommem[13336] <= 16'hFFFF;
rommem[13337] <= 16'hFFFF;
rommem[13338] <= 16'hFFFF;
rommem[13339] <= 16'hFFFF;
rommem[13340] <= 16'hFFFF;
rommem[13341] <= 16'hFFFF;
rommem[13342] <= 16'hFFFF;
rommem[13343] <= 16'hFFFF;
rommem[13344] <= 16'hFFFF;
rommem[13345] <= 16'hFFFF;
rommem[13346] <= 16'hFFFF;
rommem[13347] <= 16'hFFFF;
rommem[13348] <= 16'hFFFF;
rommem[13349] <= 16'hFFFF;
rommem[13350] <= 16'hFFFF;
rommem[13351] <= 16'hFFFF;
rommem[13352] <= 16'hFFFF;
rommem[13353] <= 16'hFFFF;
rommem[13354] <= 16'hFFFF;
rommem[13355] <= 16'hFFFF;
rommem[13356] <= 16'hFFFF;
rommem[13357] <= 16'hFFFF;
rommem[13358] <= 16'hFFFF;
rommem[13359] <= 16'hFFFF;
rommem[13360] <= 16'hFFFF;
rommem[13361] <= 16'hFFFF;
rommem[13362] <= 16'hFFFF;
rommem[13363] <= 16'hFFFF;
rommem[13364] <= 16'hFFFF;
rommem[13365] <= 16'hFFFF;
rommem[13366] <= 16'hFFFF;
rommem[13367] <= 16'hFFFF;
rommem[13368] <= 16'hFFFF;
rommem[13369] <= 16'hFFFF;
rommem[13370] <= 16'hFFFF;
rommem[13371] <= 16'hFFFF;
rommem[13372] <= 16'hFFFF;
rommem[13373] <= 16'hFFFF;
rommem[13374] <= 16'hFFFF;
rommem[13375] <= 16'hFFFF;
rommem[13376] <= 16'hFFFF;
rommem[13377] <= 16'hFFFF;
rommem[13378] <= 16'hFFFF;
rommem[13379] <= 16'hFFFF;
rommem[13380] <= 16'hFFFF;
rommem[13381] <= 16'hFFFF;
rommem[13382] <= 16'hFFFF;
rommem[13383] <= 16'hFFFF;
rommem[13384] <= 16'hFFFF;
rommem[13385] <= 16'hFFFF;
rommem[13386] <= 16'hFFFF;
rommem[13387] <= 16'hFFFF;
rommem[13388] <= 16'hFFFF;
rommem[13389] <= 16'hFFFF;
rommem[13390] <= 16'hFFFF;
rommem[13391] <= 16'hFFFF;
rommem[13392] <= 16'hFFFF;
rommem[13393] <= 16'hFFFF;
rommem[13394] <= 16'hFFFF;
rommem[13395] <= 16'hFFFF;
rommem[13396] <= 16'hFFFF;
rommem[13397] <= 16'hFFFF;
rommem[13398] <= 16'hFFFF;
rommem[13399] <= 16'hFFFF;
rommem[13400] <= 16'hFFFF;
rommem[13401] <= 16'hFFFF;
rommem[13402] <= 16'hFFFF;
rommem[13403] <= 16'hFFFF;
rommem[13404] <= 16'hFFFF;
rommem[13405] <= 16'hFFFF;
rommem[13406] <= 16'hFFFF;
rommem[13407] <= 16'hFFFF;
rommem[13408] <= 16'hFFFF;
rommem[13409] <= 16'hFFFF;
rommem[13410] <= 16'hFFFF;
rommem[13411] <= 16'hFFFF;
rommem[13412] <= 16'hFFFF;
rommem[13413] <= 16'hFFFF;
rommem[13414] <= 16'hFFFF;
rommem[13415] <= 16'hFFFF;
rommem[13416] <= 16'hFFFF;
rommem[13417] <= 16'hFFFF;
rommem[13418] <= 16'hFFFF;
rommem[13419] <= 16'hFFFF;
rommem[13420] <= 16'hFFFF;
rommem[13421] <= 16'hFFFF;
rommem[13422] <= 16'hFFFF;
rommem[13423] <= 16'hFFFF;
rommem[13424] <= 16'hFFFF;
rommem[13425] <= 16'hFFFF;
rommem[13426] <= 16'hFFFF;
rommem[13427] <= 16'hFFFF;
rommem[13428] <= 16'hFFFF;
rommem[13429] <= 16'hFFFF;
rommem[13430] <= 16'hFFFF;
rommem[13431] <= 16'hFFFF;
rommem[13432] <= 16'hFFFF;
rommem[13433] <= 16'hFFFF;
rommem[13434] <= 16'hFFFF;
rommem[13435] <= 16'hFFFF;
rommem[13436] <= 16'hFFFF;
rommem[13437] <= 16'hFFFF;
rommem[13438] <= 16'hFFFF;
rommem[13439] <= 16'hFFFF;
rommem[13440] <= 16'hFFFF;
rommem[13441] <= 16'hFFFF;
rommem[13442] <= 16'hFFFF;
rommem[13443] <= 16'hFFFF;
rommem[13444] <= 16'hFFFF;
rommem[13445] <= 16'hFFFF;
rommem[13446] <= 16'hFFFF;
rommem[13447] <= 16'hFFFF;
rommem[13448] <= 16'hFFFF;
rommem[13449] <= 16'hFFFF;
rommem[13450] <= 16'hFFFF;
rommem[13451] <= 16'hFFFF;
rommem[13452] <= 16'hFFFF;
rommem[13453] <= 16'hFFFF;
rommem[13454] <= 16'hFFFF;
rommem[13455] <= 16'hFFFF;
rommem[13456] <= 16'hFFFF;
rommem[13457] <= 16'hFFFF;
rommem[13458] <= 16'hFFFF;
rommem[13459] <= 16'hFFFF;
rommem[13460] <= 16'hFFFF;
rommem[13461] <= 16'hFFFF;
rommem[13462] <= 16'hFFFF;
rommem[13463] <= 16'hFFFF;
rommem[13464] <= 16'hFFFF;
rommem[13465] <= 16'hFFFF;
rommem[13466] <= 16'hFFFF;
rommem[13467] <= 16'hFFFF;
rommem[13468] <= 16'hFFFF;
rommem[13469] <= 16'hFFFF;
rommem[13470] <= 16'hFFFF;
rommem[13471] <= 16'hFFFF;
rommem[13472] <= 16'hFFFF;
rommem[13473] <= 16'hFFFF;
rommem[13474] <= 16'hFFFF;
rommem[13475] <= 16'hFFFF;
rommem[13476] <= 16'hFFFF;
rommem[13477] <= 16'hFFFF;
rommem[13478] <= 16'hFFFF;
rommem[13479] <= 16'hFFFF;
rommem[13480] <= 16'hFFFF;
rommem[13481] <= 16'hFFFF;
rommem[13482] <= 16'hFFFF;
rommem[13483] <= 16'hFFFF;
rommem[13484] <= 16'hFFFF;
rommem[13485] <= 16'hFFFF;
rommem[13486] <= 16'hFFFF;
rommem[13487] <= 16'hFFFF;
rommem[13488] <= 16'hFFFF;
rommem[13489] <= 16'hFFFF;
rommem[13490] <= 16'hFFFF;
rommem[13491] <= 16'hFFFF;
rommem[13492] <= 16'hFFFF;
rommem[13493] <= 16'hFFFF;
rommem[13494] <= 16'hFFFF;
rommem[13495] <= 16'hFFFF;
rommem[13496] <= 16'hFFFF;
rommem[13497] <= 16'hFFFF;
rommem[13498] <= 16'hFFFF;
rommem[13499] <= 16'hFFFF;
rommem[13500] <= 16'hFFFF;
rommem[13501] <= 16'hFFFF;
rommem[13502] <= 16'hFFFF;
rommem[13503] <= 16'hFFFF;
rommem[13504] <= 16'hFFFF;
rommem[13505] <= 16'hFFFF;
rommem[13506] <= 16'hFFFF;
rommem[13507] <= 16'hFFFF;
rommem[13508] <= 16'hFFFF;
rommem[13509] <= 16'hFFFF;
rommem[13510] <= 16'hFFFF;
rommem[13511] <= 16'hFFFF;
rommem[13512] <= 16'hFFFF;
rommem[13513] <= 16'hFFFF;
rommem[13514] <= 16'hFFFF;
rommem[13515] <= 16'hFFFF;
rommem[13516] <= 16'hFFFF;
rommem[13517] <= 16'hFFFF;
rommem[13518] <= 16'hFFFF;
rommem[13519] <= 16'hFFFF;
rommem[13520] <= 16'hFFFF;
rommem[13521] <= 16'hFFFF;
rommem[13522] <= 16'hFFFF;
rommem[13523] <= 16'hFFFF;
rommem[13524] <= 16'hFFFF;
rommem[13525] <= 16'hFFFF;
rommem[13526] <= 16'hFFFF;
rommem[13527] <= 16'hFFFF;
rommem[13528] <= 16'hFFFF;
rommem[13529] <= 16'hFFFF;
rommem[13530] <= 16'hFFFF;
rommem[13531] <= 16'hFFFF;
rommem[13532] <= 16'hFFFF;
rommem[13533] <= 16'hFFFF;
rommem[13534] <= 16'hFFFF;
rommem[13535] <= 16'hFFFF;
rommem[13536] <= 16'hFFFF;
rommem[13537] <= 16'hFFFF;
rommem[13538] <= 16'hFFFF;
rommem[13539] <= 16'hFFFF;
rommem[13540] <= 16'hFFFF;
rommem[13541] <= 16'hFFFF;
rommem[13542] <= 16'hFFFF;
rommem[13543] <= 16'hFFFF;
rommem[13544] <= 16'hFFFF;
rommem[13545] <= 16'hFFFF;
rommem[13546] <= 16'hFFFF;
rommem[13547] <= 16'hFFFF;
rommem[13548] <= 16'hFFFF;
rommem[13549] <= 16'hFFFF;
rommem[13550] <= 16'hFFFF;
rommem[13551] <= 16'hFFFF;
rommem[13552] <= 16'hFFFF;
rommem[13553] <= 16'hFFFF;
rommem[13554] <= 16'hFFFF;
rommem[13555] <= 16'hFFFF;
rommem[13556] <= 16'hFFFF;
rommem[13557] <= 16'hFFFF;
rommem[13558] <= 16'hFFFF;
rommem[13559] <= 16'hFFFF;
rommem[13560] <= 16'hFFFF;
rommem[13561] <= 16'hFFFF;
rommem[13562] <= 16'hFFFF;
rommem[13563] <= 16'hFFFF;
rommem[13564] <= 16'hFFFF;
rommem[13565] <= 16'hFFFF;
rommem[13566] <= 16'hFFFF;
rommem[13567] <= 16'hFFFF;
rommem[13568] <= 16'hFFFF;
rommem[13569] <= 16'hFFFF;
rommem[13570] <= 16'hFFFF;
rommem[13571] <= 16'hFFFF;
rommem[13572] <= 16'hFFFF;
rommem[13573] <= 16'hFFFF;
rommem[13574] <= 16'hFFFF;
rommem[13575] <= 16'hFFFF;
rommem[13576] <= 16'hFFFF;
rommem[13577] <= 16'hFFFF;
rommem[13578] <= 16'hFFFF;
rommem[13579] <= 16'hFFFF;
rommem[13580] <= 16'hFFFF;
rommem[13581] <= 16'hFFFF;
rommem[13582] <= 16'hFFFF;
rommem[13583] <= 16'hFFFF;
rommem[13584] <= 16'hFFFF;
rommem[13585] <= 16'hFFFF;
rommem[13586] <= 16'hFFFF;
rommem[13587] <= 16'hFFFF;
rommem[13588] <= 16'hFFFF;
rommem[13589] <= 16'hFFFF;
rommem[13590] <= 16'hFFFF;
rommem[13591] <= 16'hFFFF;
rommem[13592] <= 16'hFFFF;
rommem[13593] <= 16'hFFFF;
rommem[13594] <= 16'hFFFF;
rommem[13595] <= 16'hFFFF;
rommem[13596] <= 16'hFFFF;
rommem[13597] <= 16'hFFFF;
rommem[13598] <= 16'hFFFF;
rommem[13599] <= 16'hFFFF;
rommem[13600] <= 16'hFFFF;
rommem[13601] <= 16'hFFFF;
rommem[13602] <= 16'hFFFF;
rommem[13603] <= 16'hFFFF;
rommem[13604] <= 16'hFFFF;
rommem[13605] <= 16'hFFFF;
rommem[13606] <= 16'hFFFF;
rommem[13607] <= 16'hFFFF;
rommem[13608] <= 16'hFFFF;
rommem[13609] <= 16'hFFFF;
rommem[13610] <= 16'hFFFF;
rommem[13611] <= 16'hFFFF;
rommem[13612] <= 16'hFFFF;
rommem[13613] <= 16'hFFFF;
rommem[13614] <= 16'hFFFF;
rommem[13615] <= 16'hFFFF;
rommem[13616] <= 16'hFFFF;
rommem[13617] <= 16'hFFFF;
rommem[13618] <= 16'hFFFF;
rommem[13619] <= 16'hFFFF;
rommem[13620] <= 16'hFFFF;
rommem[13621] <= 16'hFFFF;
rommem[13622] <= 16'hFFFF;
rommem[13623] <= 16'hFFFF;
rommem[13624] <= 16'hFFFF;
rommem[13625] <= 16'hFFFF;
rommem[13626] <= 16'hFFFF;
rommem[13627] <= 16'hFFFF;
rommem[13628] <= 16'hFFFF;
rommem[13629] <= 16'hFFFF;
rommem[13630] <= 16'hFFFF;
rommem[13631] <= 16'hFFFF;
rommem[13632] <= 16'hFFFF;
rommem[13633] <= 16'hFFFF;
rommem[13634] <= 16'hFFFF;
rommem[13635] <= 16'hFFFF;
rommem[13636] <= 16'hFFFF;
rommem[13637] <= 16'hFFFF;
rommem[13638] <= 16'hFFFF;
rommem[13639] <= 16'hFFFF;
rommem[13640] <= 16'hFFFF;
rommem[13641] <= 16'hFFFF;
rommem[13642] <= 16'hFFFF;
rommem[13643] <= 16'hFFFF;
rommem[13644] <= 16'hFFFF;
rommem[13645] <= 16'hFFFF;
rommem[13646] <= 16'hFFFF;
rommem[13647] <= 16'hFFFF;
rommem[13648] <= 16'hFFFF;
rommem[13649] <= 16'hFFFF;
rommem[13650] <= 16'hFFFF;
rommem[13651] <= 16'hFFFF;
rommem[13652] <= 16'hFFFF;
rommem[13653] <= 16'hFFFF;
rommem[13654] <= 16'hFFFF;
rommem[13655] <= 16'hFFFF;
rommem[13656] <= 16'hFFFF;
rommem[13657] <= 16'hFFFF;
rommem[13658] <= 16'hFFFF;
rommem[13659] <= 16'hFFFF;
rommem[13660] <= 16'hFFFF;
rommem[13661] <= 16'hFFFF;
rommem[13662] <= 16'hFFFF;
rommem[13663] <= 16'hFFFF;
rommem[13664] <= 16'hFFFF;
rommem[13665] <= 16'hFFFF;
rommem[13666] <= 16'hFFFF;
rommem[13667] <= 16'hFFFF;
rommem[13668] <= 16'hFFFF;
rommem[13669] <= 16'hFFFF;
rommem[13670] <= 16'hFFFF;
rommem[13671] <= 16'hFFFF;
rommem[13672] <= 16'hFFFF;
rommem[13673] <= 16'hFFFF;
rommem[13674] <= 16'hFFFF;
rommem[13675] <= 16'hFFFF;
rommem[13676] <= 16'hFFFF;
rommem[13677] <= 16'hFFFF;
rommem[13678] <= 16'hFFFF;
rommem[13679] <= 16'hFFFF;
rommem[13680] <= 16'hFFFF;
rommem[13681] <= 16'hFFFF;
rommem[13682] <= 16'hFFFF;
rommem[13683] <= 16'hFFFF;
rommem[13684] <= 16'hFFFF;
rommem[13685] <= 16'hFFFF;
rommem[13686] <= 16'hFFFF;
rommem[13687] <= 16'hFFFF;
rommem[13688] <= 16'hFFFF;
rommem[13689] <= 16'hFFFF;
rommem[13690] <= 16'hFFFF;
rommem[13691] <= 16'hFFFF;
rommem[13692] <= 16'hFFFF;
rommem[13693] <= 16'hFFFF;
rommem[13694] <= 16'hFFFF;
rommem[13695] <= 16'hFFFF;
rommem[13696] <= 16'hFFFF;
rommem[13697] <= 16'hFFFF;
rommem[13698] <= 16'hFFFF;
rommem[13699] <= 16'hFFFF;
rommem[13700] <= 16'hFFFF;
rommem[13701] <= 16'hFFFF;
rommem[13702] <= 16'hFFFF;
rommem[13703] <= 16'hFFFF;
rommem[13704] <= 16'hFFFF;
rommem[13705] <= 16'hFFFF;
rommem[13706] <= 16'hFFFF;
rommem[13707] <= 16'hFFFF;
rommem[13708] <= 16'hFFFF;
rommem[13709] <= 16'hFFFF;
rommem[13710] <= 16'hFFFF;
rommem[13711] <= 16'hFFFF;
rommem[13712] <= 16'hFFFF;
rommem[13713] <= 16'hFFFF;
rommem[13714] <= 16'hFFFF;
rommem[13715] <= 16'hFFFF;
rommem[13716] <= 16'hFFFF;
rommem[13717] <= 16'hFFFF;
rommem[13718] <= 16'hFFFF;
rommem[13719] <= 16'hFFFF;
rommem[13720] <= 16'hFFFF;
rommem[13721] <= 16'hFFFF;
rommem[13722] <= 16'hFFFF;
rommem[13723] <= 16'hFFFF;
rommem[13724] <= 16'hFFFF;
rommem[13725] <= 16'hFFFF;
rommem[13726] <= 16'hFFFF;
rommem[13727] <= 16'hFFFF;
rommem[13728] <= 16'hFFFF;
rommem[13729] <= 16'hFFFF;
rommem[13730] <= 16'hFFFF;
rommem[13731] <= 16'hFFFF;
rommem[13732] <= 16'hFFFF;
rommem[13733] <= 16'hFFFF;
rommem[13734] <= 16'hFFFF;
rommem[13735] <= 16'hFFFF;
rommem[13736] <= 16'hFFFF;
rommem[13737] <= 16'hFFFF;
rommem[13738] <= 16'hFFFF;
rommem[13739] <= 16'hFFFF;
rommem[13740] <= 16'hFFFF;
rommem[13741] <= 16'hFFFF;
rommem[13742] <= 16'hFFFF;
rommem[13743] <= 16'hFFFF;
rommem[13744] <= 16'hFFFF;
rommem[13745] <= 16'hFFFF;
rommem[13746] <= 16'hFFFF;
rommem[13747] <= 16'hFFFF;
rommem[13748] <= 16'hFFFF;
rommem[13749] <= 16'hFFFF;
rommem[13750] <= 16'hFFFF;
rommem[13751] <= 16'hFFFF;
rommem[13752] <= 16'hFFFF;
rommem[13753] <= 16'hFFFF;
rommem[13754] <= 16'hFFFF;
rommem[13755] <= 16'hFFFF;
rommem[13756] <= 16'hFFFF;
rommem[13757] <= 16'hFFFF;
rommem[13758] <= 16'hFFFF;
rommem[13759] <= 16'hFFFF;
rommem[13760] <= 16'hFFFF;
rommem[13761] <= 16'hFFFF;
rommem[13762] <= 16'hFFFF;
rommem[13763] <= 16'hFFFF;
rommem[13764] <= 16'hFFFF;
rommem[13765] <= 16'hFFFF;
rommem[13766] <= 16'hFFFF;
rommem[13767] <= 16'hFFFF;
rommem[13768] <= 16'hFFFF;
rommem[13769] <= 16'hFFFF;
rommem[13770] <= 16'hFFFF;
rommem[13771] <= 16'hFFFF;
rommem[13772] <= 16'hFFFF;
rommem[13773] <= 16'hFFFF;
rommem[13774] <= 16'hFFFF;
rommem[13775] <= 16'hFFFF;
rommem[13776] <= 16'hFFFF;
rommem[13777] <= 16'hFFFF;
rommem[13778] <= 16'hFFFF;
rommem[13779] <= 16'hFFFF;
rommem[13780] <= 16'hFFFF;
rommem[13781] <= 16'hFFFF;
rommem[13782] <= 16'hFFFF;
rommem[13783] <= 16'hFFFF;
rommem[13784] <= 16'hFFFF;
rommem[13785] <= 16'hFFFF;
rommem[13786] <= 16'hFFFF;
rommem[13787] <= 16'hFFFF;
rommem[13788] <= 16'hFFFF;
rommem[13789] <= 16'hFFFF;
rommem[13790] <= 16'hFFFF;
rommem[13791] <= 16'hFFFF;
rommem[13792] <= 16'hFFFF;
rommem[13793] <= 16'hFFFF;
rommem[13794] <= 16'hFFFF;
rommem[13795] <= 16'hFFFF;
rommem[13796] <= 16'hFFFF;
rommem[13797] <= 16'hFFFF;
rommem[13798] <= 16'hFFFF;
rommem[13799] <= 16'hFFFF;
rommem[13800] <= 16'hFFFF;
rommem[13801] <= 16'hFFFF;
rommem[13802] <= 16'hFFFF;
rommem[13803] <= 16'hFFFF;
rommem[13804] <= 16'hFFFF;
rommem[13805] <= 16'hFFFF;
rommem[13806] <= 16'hFFFF;
rommem[13807] <= 16'hFFFF;
rommem[13808] <= 16'hFFFF;
rommem[13809] <= 16'hFFFF;
rommem[13810] <= 16'hFFFF;
rommem[13811] <= 16'hFFFF;
rommem[13812] <= 16'hFFFF;
rommem[13813] <= 16'hFFFF;
rommem[13814] <= 16'hFFFF;
rommem[13815] <= 16'hFFFF;
rommem[13816] <= 16'hFFFF;
rommem[13817] <= 16'hFFFF;
rommem[13818] <= 16'hFFFF;
rommem[13819] <= 16'hFFFF;
rommem[13820] <= 16'hFFFF;
rommem[13821] <= 16'hFFFF;
rommem[13822] <= 16'hFFFF;
rommem[13823] <= 16'hFFFF;
rommem[13824] <= 16'hFFFF;
rommem[13825] <= 16'hFFFF;
rommem[13826] <= 16'hFFFF;
rommem[13827] <= 16'hFFFF;
rommem[13828] <= 16'hFFFF;
rommem[13829] <= 16'hFFFF;
rommem[13830] <= 16'hFFFF;
rommem[13831] <= 16'hFFFF;
rommem[13832] <= 16'hFFFF;
rommem[13833] <= 16'hFFFF;
rommem[13834] <= 16'hFFFF;
rommem[13835] <= 16'hFFFF;
rommem[13836] <= 16'hFFFF;
rommem[13837] <= 16'hFFFF;
rommem[13838] <= 16'hFFFF;
rommem[13839] <= 16'hFFFF;
rommem[13840] <= 16'hFFFF;
rommem[13841] <= 16'hFFFF;
rommem[13842] <= 16'hFFFF;
rommem[13843] <= 16'hFFFF;
rommem[13844] <= 16'hFFFF;
rommem[13845] <= 16'hFFFF;
rommem[13846] <= 16'hFFFF;
rommem[13847] <= 16'hFFFF;
rommem[13848] <= 16'hFFFF;
rommem[13849] <= 16'hFFFF;
rommem[13850] <= 16'hFFFF;
rommem[13851] <= 16'hFFFF;
rommem[13852] <= 16'hFFFF;
rommem[13853] <= 16'hFFFF;
rommem[13854] <= 16'hFFFF;
rommem[13855] <= 16'hFFFF;
rommem[13856] <= 16'hFFFF;
rommem[13857] <= 16'hFFFF;
rommem[13858] <= 16'hFFFF;
rommem[13859] <= 16'hFFFF;
rommem[13860] <= 16'hFFFF;
rommem[13861] <= 16'hFFFF;
rommem[13862] <= 16'hFFFF;
rommem[13863] <= 16'hFFFF;
rommem[13864] <= 16'hFFFF;
rommem[13865] <= 16'hFFFF;
rommem[13866] <= 16'hFFFF;
rommem[13867] <= 16'hFFFF;
rommem[13868] <= 16'hFFFF;
rommem[13869] <= 16'hFFFF;
rommem[13870] <= 16'hFFFF;
rommem[13871] <= 16'hFFFF;
rommem[13872] <= 16'hFFFF;
rommem[13873] <= 16'hFFFF;
rommem[13874] <= 16'hFFFF;
rommem[13875] <= 16'hFFFF;
rommem[13876] <= 16'hFFFF;
rommem[13877] <= 16'hFFFF;
rommem[13878] <= 16'hFFFF;
rommem[13879] <= 16'hFFFF;
rommem[13880] <= 16'hFFFF;
rommem[13881] <= 16'hFFFF;
rommem[13882] <= 16'hFFFF;
rommem[13883] <= 16'hFFFF;
rommem[13884] <= 16'hFFFF;
rommem[13885] <= 16'hFFFF;
rommem[13886] <= 16'hFFFF;
rommem[13887] <= 16'hFFFF;
rommem[13888] <= 16'hFFFF;
rommem[13889] <= 16'hFFFF;
rommem[13890] <= 16'hFFFF;
rommem[13891] <= 16'hFFFF;
rommem[13892] <= 16'hFFFF;
rommem[13893] <= 16'hFFFF;
rommem[13894] <= 16'hFFFF;
rommem[13895] <= 16'hFFFF;
rommem[13896] <= 16'hFFFF;
rommem[13897] <= 16'hFFFF;
rommem[13898] <= 16'hFFFF;
rommem[13899] <= 16'hFFFF;
rommem[13900] <= 16'hFFFF;
rommem[13901] <= 16'hFFFF;
rommem[13902] <= 16'hFFFF;
rommem[13903] <= 16'hFFFF;
rommem[13904] <= 16'hFFFF;
rommem[13905] <= 16'hFFFF;
rommem[13906] <= 16'hFFFF;
rommem[13907] <= 16'hFFFF;
rommem[13908] <= 16'hFFFF;
rommem[13909] <= 16'hFFFF;
rommem[13910] <= 16'hFFFF;
rommem[13911] <= 16'hFFFF;
rommem[13912] <= 16'hFFFF;
rommem[13913] <= 16'hFFFF;
rommem[13914] <= 16'hFFFF;
rommem[13915] <= 16'hFFFF;
rommem[13916] <= 16'hFFFF;
rommem[13917] <= 16'hFFFF;
rommem[13918] <= 16'hFFFF;
rommem[13919] <= 16'hFFFF;
rommem[13920] <= 16'hFFFF;
rommem[13921] <= 16'hFFFF;
rommem[13922] <= 16'hFFFF;
rommem[13923] <= 16'hFFFF;
rommem[13924] <= 16'hFFFF;
rommem[13925] <= 16'hFFFF;
rommem[13926] <= 16'hFFFF;
rommem[13927] <= 16'hFFFF;
rommem[13928] <= 16'hFFFF;
rommem[13929] <= 16'hFFFF;
rommem[13930] <= 16'hFFFF;
rommem[13931] <= 16'hFFFF;
rommem[13932] <= 16'hFFFF;
rommem[13933] <= 16'hFFFF;
rommem[13934] <= 16'hFFFF;
rommem[13935] <= 16'hFFFF;
rommem[13936] <= 16'hFFFF;
rommem[13937] <= 16'hFFFF;
rommem[13938] <= 16'hFFFF;
rommem[13939] <= 16'hFFFF;
rommem[13940] <= 16'hFFFF;
rommem[13941] <= 16'hFFFF;
rommem[13942] <= 16'hFFFF;
rommem[13943] <= 16'hFFFF;
rommem[13944] <= 16'hFFFF;
rommem[13945] <= 16'hFFFF;
rommem[13946] <= 16'hFFFF;
rommem[13947] <= 16'hFFFF;
rommem[13948] <= 16'hFFFF;
rommem[13949] <= 16'hFFFF;
rommem[13950] <= 16'hFFFF;
rommem[13951] <= 16'hFFFF;
rommem[13952] <= 16'hFFFF;
rommem[13953] <= 16'hFFFF;
rommem[13954] <= 16'hFFFF;
rommem[13955] <= 16'hFFFF;
rommem[13956] <= 16'hFFFF;
rommem[13957] <= 16'hFFFF;
rommem[13958] <= 16'hFFFF;
rommem[13959] <= 16'hFFFF;
rommem[13960] <= 16'hFFFF;
rommem[13961] <= 16'hFFFF;
rommem[13962] <= 16'hFFFF;
rommem[13963] <= 16'hFFFF;
rommem[13964] <= 16'hFFFF;
rommem[13965] <= 16'hFFFF;
rommem[13966] <= 16'hFFFF;
rommem[13967] <= 16'hFFFF;
rommem[13968] <= 16'hFFFF;
rommem[13969] <= 16'hFFFF;
rommem[13970] <= 16'hFFFF;
rommem[13971] <= 16'hFFFF;
rommem[13972] <= 16'hFFFF;
rommem[13973] <= 16'hFFFF;
rommem[13974] <= 16'hFFFF;
rommem[13975] <= 16'hFFFF;
rommem[13976] <= 16'hFFFF;
rommem[13977] <= 16'hFFFF;
rommem[13978] <= 16'hFFFF;
rommem[13979] <= 16'hFFFF;
rommem[13980] <= 16'hFFFF;
rommem[13981] <= 16'hFFFF;
rommem[13982] <= 16'hFFFF;
rommem[13983] <= 16'hFFFF;
rommem[13984] <= 16'hFFFF;
rommem[13985] <= 16'hFFFF;
rommem[13986] <= 16'hFFFF;
rommem[13987] <= 16'hFFFF;
rommem[13988] <= 16'hFFFF;
rommem[13989] <= 16'hFFFF;
rommem[13990] <= 16'hFFFF;
rommem[13991] <= 16'hFFFF;
rommem[13992] <= 16'hFFFF;
rommem[13993] <= 16'hFFFF;
rommem[13994] <= 16'hFFFF;
rommem[13995] <= 16'hFFFF;
rommem[13996] <= 16'hFFFF;
rommem[13997] <= 16'hFFFF;
rommem[13998] <= 16'hFFFF;
rommem[13999] <= 16'hFFFF;
rommem[14000] <= 16'hFFFF;
rommem[14001] <= 16'hFFFF;
rommem[14002] <= 16'hFFFF;
rommem[14003] <= 16'hFFFF;
rommem[14004] <= 16'hFFFF;
rommem[14005] <= 16'hFFFF;
rommem[14006] <= 16'hFFFF;
rommem[14007] <= 16'hFFFF;
rommem[14008] <= 16'hFFFF;
rommem[14009] <= 16'hFFFF;
rommem[14010] <= 16'hFFFF;
rommem[14011] <= 16'hFFFF;
rommem[14012] <= 16'hFFFF;
rommem[14013] <= 16'hFFFF;
rommem[14014] <= 16'hFFFF;
rommem[14015] <= 16'hFFFF;
rommem[14016] <= 16'hFFFF;
rommem[14017] <= 16'hFFFF;
rommem[14018] <= 16'hFFFF;
rommem[14019] <= 16'hFFFF;
rommem[14020] <= 16'hFFFF;
rommem[14021] <= 16'hFFFF;
rommem[14022] <= 16'hFFFF;
rommem[14023] <= 16'hFFFF;
rommem[14024] <= 16'hFFFF;
rommem[14025] <= 16'hFFFF;
rommem[14026] <= 16'hFFFF;
rommem[14027] <= 16'hFFFF;
rommem[14028] <= 16'hFFFF;
rommem[14029] <= 16'hFFFF;
rommem[14030] <= 16'hFFFF;
rommem[14031] <= 16'hFFFF;
rommem[14032] <= 16'hFFFF;
rommem[14033] <= 16'hFFFF;
rommem[14034] <= 16'hFFFF;
rommem[14035] <= 16'hFFFF;
rommem[14036] <= 16'hFFFF;
rommem[14037] <= 16'hFFFF;
rommem[14038] <= 16'hFFFF;
rommem[14039] <= 16'hFFFF;
rommem[14040] <= 16'hFFFF;
rommem[14041] <= 16'hFFFF;
rommem[14042] <= 16'hFFFF;
rommem[14043] <= 16'hFFFF;
rommem[14044] <= 16'hFFFF;
rommem[14045] <= 16'hFFFF;
rommem[14046] <= 16'hFFFF;
rommem[14047] <= 16'hFFFF;
rommem[14048] <= 16'hFFFF;
rommem[14049] <= 16'hFFFF;
rommem[14050] <= 16'hFFFF;
rommem[14051] <= 16'hFFFF;
rommem[14052] <= 16'hFFFF;
rommem[14053] <= 16'hFFFF;
rommem[14054] <= 16'hFFFF;
rommem[14055] <= 16'hFFFF;
rommem[14056] <= 16'hFFFF;
rommem[14057] <= 16'hFFFF;
rommem[14058] <= 16'hFFFF;
rommem[14059] <= 16'hFFFF;
rommem[14060] <= 16'hFFFF;
rommem[14061] <= 16'hFFFF;
rommem[14062] <= 16'hFFFF;
rommem[14063] <= 16'hFFFF;
rommem[14064] <= 16'hFFFF;
rommem[14065] <= 16'hFFFF;
rommem[14066] <= 16'hFFFF;
rommem[14067] <= 16'hFFFF;
rommem[14068] <= 16'hFFFF;
rommem[14069] <= 16'hFFFF;
rommem[14070] <= 16'hFFFF;
rommem[14071] <= 16'hFFFF;
rommem[14072] <= 16'hFFFF;
rommem[14073] <= 16'hFFFF;
rommem[14074] <= 16'hFFFF;
rommem[14075] <= 16'hFFFF;
rommem[14076] <= 16'hFFFF;
rommem[14077] <= 16'hFFFF;
rommem[14078] <= 16'hFFFF;
rommem[14079] <= 16'hFFFF;
rommem[14080] <= 16'hFFFF;
rommem[14081] <= 16'hFFFF;
rommem[14082] <= 16'hFFFF;
rommem[14083] <= 16'hFFFF;
rommem[14084] <= 16'hFFFF;
rommem[14085] <= 16'hFFFF;
rommem[14086] <= 16'hFFFF;
rommem[14087] <= 16'hFFFF;
rommem[14088] <= 16'hFFFF;
rommem[14089] <= 16'hFFFF;
rommem[14090] <= 16'hFFFF;
rommem[14091] <= 16'hFFFF;
rommem[14092] <= 16'hFFFF;
rommem[14093] <= 16'hFFFF;
rommem[14094] <= 16'hFFFF;
rommem[14095] <= 16'hFFFF;
rommem[14096] <= 16'hFFFF;
rommem[14097] <= 16'hFFFF;
rommem[14098] <= 16'hFFFF;
rommem[14099] <= 16'hFFFF;
rommem[14100] <= 16'hFFFF;
rommem[14101] <= 16'hFFFF;
rommem[14102] <= 16'hFFFF;
rommem[14103] <= 16'hFFFF;
rommem[14104] <= 16'hFFFF;
rommem[14105] <= 16'hFFFF;
rommem[14106] <= 16'hFFFF;
rommem[14107] <= 16'hFFFF;
rommem[14108] <= 16'hFFFF;
rommem[14109] <= 16'hFFFF;
rommem[14110] <= 16'hFFFF;
rommem[14111] <= 16'hFFFF;
rommem[14112] <= 16'hFFFF;
rommem[14113] <= 16'hFFFF;
rommem[14114] <= 16'hFFFF;
rommem[14115] <= 16'hFFFF;
rommem[14116] <= 16'hFFFF;
rommem[14117] <= 16'hFFFF;
rommem[14118] <= 16'hFFFF;
rommem[14119] <= 16'hFFFF;
rommem[14120] <= 16'hFFFF;
rommem[14121] <= 16'hFFFF;
rommem[14122] <= 16'hFFFF;
rommem[14123] <= 16'hFFFF;
rommem[14124] <= 16'hFFFF;
rommem[14125] <= 16'hFFFF;
rommem[14126] <= 16'hFFFF;
rommem[14127] <= 16'hFFFF;
rommem[14128] <= 16'hFFFF;
rommem[14129] <= 16'hFFFF;
rommem[14130] <= 16'hFFFF;
rommem[14131] <= 16'hFFFF;
rommem[14132] <= 16'hFFFF;
rommem[14133] <= 16'hFFFF;
rommem[14134] <= 16'hFFFF;
rommem[14135] <= 16'hFFFF;
rommem[14136] <= 16'hFFFF;
rommem[14137] <= 16'hFFFF;
rommem[14138] <= 16'hFFFF;
rommem[14139] <= 16'hFFFF;
rommem[14140] <= 16'hFFFF;
rommem[14141] <= 16'hFFFF;
rommem[14142] <= 16'hFFFF;
rommem[14143] <= 16'hFFFF;
rommem[14144] <= 16'hFFFF;
rommem[14145] <= 16'hFFFF;
rommem[14146] <= 16'hFFFF;
rommem[14147] <= 16'hFFFF;
rommem[14148] <= 16'hFFFF;
rommem[14149] <= 16'hFFFF;
rommem[14150] <= 16'hFFFF;
rommem[14151] <= 16'hFFFF;
rommem[14152] <= 16'hFFFF;
rommem[14153] <= 16'hFFFF;
rommem[14154] <= 16'hFFFF;
rommem[14155] <= 16'hFFFF;
rommem[14156] <= 16'hFFFF;
rommem[14157] <= 16'hFFFF;
rommem[14158] <= 16'hFFFF;
rommem[14159] <= 16'hFFFF;
rommem[14160] <= 16'hFFFF;
rommem[14161] <= 16'hFFFF;
rommem[14162] <= 16'hFFFF;
rommem[14163] <= 16'hFFFF;
rommem[14164] <= 16'hFFFF;
rommem[14165] <= 16'hFFFF;
rommem[14166] <= 16'hFFFF;
rommem[14167] <= 16'hFFFF;
rommem[14168] <= 16'hFFFF;
rommem[14169] <= 16'hFFFF;
rommem[14170] <= 16'hFFFF;
rommem[14171] <= 16'hFFFF;
rommem[14172] <= 16'hFFFF;
rommem[14173] <= 16'hFFFF;
rommem[14174] <= 16'hFFFF;
rommem[14175] <= 16'hFFFF;
rommem[14176] <= 16'hFFFF;
rommem[14177] <= 16'hFFFF;
rommem[14178] <= 16'hFFFF;
rommem[14179] <= 16'hFFFF;
rommem[14180] <= 16'hFFFF;
rommem[14181] <= 16'hFFFF;
rommem[14182] <= 16'hFFFF;
rommem[14183] <= 16'hFFFF;
rommem[14184] <= 16'hFFFF;
rommem[14185] <= 16'hFFFF;
rommem[14186] <= 16'hFFFF;
rommem[14187] <= 16'hFFFF;
rommem[14188] <= 16'hFFFF;
rommem[14189] <= 16'hFFFF;
rommem[14190] <= 16'hFFFF;
rommem[14191] <= 16'hFFFF;
rommem[14192] <= 16'hFFFF;
rommem[14193] <= 16'hFFFF;
rommem[14194] <= 16'hFFFF;
rommem[14195] <= 16'hFFFF;
rommem[14196] <= 16'hFFFF;
rommem[14197] <= 16'hFFFF;
rommem[14198] <= 16'hFFFF;
rommem[14199] <= 16'hFFFF;
rommem[14200] <= 16'hFFFF;
rommem[14201] <= 16'hFFFF;
rommem[14202] <= 16'hFFFF;
rommem[14203] <= 16'hFFFF;
rommem[14204] <= 16'hFFFF;
rommem[14205] <= 16'hFFFF;
rommem[14206] <= 16'hFFFF;
rommem[14207] <= 16'hFFFF;
rommem[14208] <= 16'hFFFF;
rommem[14209] <= 16'hFFFF;
rommem[14210] <= 16'hFFFF;
rommem[14211] <= 16'hFFFF;
rommem[14212] <= 16'hFFFF;
rommem[14213] <= 16'hFFFF;
rommem[14214] <= 16'hFFFF;
rommem[14215] <= 16'hFFFF;
rommem[14216] <= 16'hFFFF;
rommem[14217] <= 16'hFFFF;
rommem[14218] <= 16'hFFFF;
rommem[14219] <= 16'hFFFF;
rommem[14220] <= 16'hFFFF;
rommem[14221] <= 16'hFFFF;
rommem[14222] <= 16'hFFFF;
rommem[14223] <= 16'hFFFF;
rommem[14224] <= 16'hFFFF;
rommem[14225] <= 16'hFFFF;
rommem[14226] <= 16'hFFFF;
rommem[14227] <= 16'hFFFF;
rommem[14228] <= 16'hFFFF;
rommem[14229] <= 16'hFFFF;
rommem[14230] <= 16'hFFFF;
rommem[14231] <= 16'hFFFF;
rommem[14232] <= 16'hFFFF;
rommem[14233] <= 16'hFFFF;
rommem[14234] <= 16'hFFFF;
rommem[14235] <= 16'hFFFF;
rommem[14236] <= 16'hFFFF;
rommem[14237] <= 16'hFFFF;
rommem[14238] <= 16'hFFFF;
rommem[14239] <= 16'hFFFF;
rommem[14240] <= 16'hFFFF;
rommem[14241] <= 16'hFFFF;
rommem[14242] <= 16'hFFFF;
rommem[14243] <= 16'hFFFF;
rommem[14244] <= 16'hFFFF;
rommem[14245] <= 16'hFFFF;
rommem[14246] <= 16'hFFFF;
rommem[14247] <= 16'hFFFF;
rommem[14248] <= 16'hFFFF;
rommem[14249] <= 16'hFFFF;
rommem[14250] <= 16'hFFFF;
rommem[14251] <= 16'hFFFF;
rommem[14252] <= 16'hFFFF;
rommem[14253] <= 16'hFFFF;
rommem[14254] <= 16'hFFFF;
rommem[14255] <= 16'hFFFF;
rommem[14256] <= 16'hFFFF;
rommem[14257] <= 16'hFFFF;
rommem[14258] <= 16'hFFFF;
rommem[14259] <= 16'hFFFF;
rommem[14260] <= 16'hFFFF;
rommem[14261] <= 16'hFFFF;
rommem[14262] <= 16'hFFFF;
rommem[14263] <= 16'hFFFF;
rommem[14264] <= 16'hFFFF;
rommem[14265] <= 16'hFFFF;
rommem[14266] <= 16'hFFFF;
rommem[14267] <= 16'hFFFF;
rommem[14268] <= 16'hFFFF;
rommem[14269] <= 16'hFFFF;
rommem[14270] <= 16'hFFFF;
rommem[14271] <= 16'hFFFF;
rommem[14272] <= 16'hFFFF;
rommem[14273] <= 16'hFFFF;
rommem[14274] <= 16'hFFFF;
rommem[14275] <= 16'hFFFF;
rommem[14276] <= 16'hFFFF;
rommem[14277] <= 16'hFFFF;
rommem[14278] <= 16'hFFFF;
rommem[14279] <= 16'hFFFF;
rommem[14280] <= 16'hFFFF;
rommem[14281] <= 16'hFFFF;
rommem[14282] <= 16'hFFFF;
rommem[14283] <= 16'hFFFF;
rommem[14284] <= 16'hFFFF;
rommem[14285] <= 16'hFFFF;
rommem[14286] <= 16'hFFFF;
rommem[14287] <= 16'hFFFF;
rommem[14288] <= 16'hFFFF;
rommem[14289] <= 16'hFFFF;
rommem[14290] <= 16'hFFFF;
rommem[14291] <= 16'hFFFF;
rommem[14292] <= 16'hFFFF;
rommem[14293] <= 16'hFFFF;
rommem[14294] <= 16'hFFFF;
rommem[14295] <= 16'hFFFF;
rommem[14296] <= 16'hFFFF;
rommem[14297] <= 16'hFFFF;
rommem[14298] <= 16'hFFFF;
rommem[14299] <= 16'hFFFF;
rommem[14300] <= 16'hFFFF;
rommem[14301] <= 16'hFFFF;
rommem[14302] <= 16'hFFFF;
rommem[14303] <= 16'hFFFF;
rommem[14304] <= 16'hFFFF;
rommem[14305] <= 16'hFFFF;
rommem[14306] <= 16'hFFFF;
rommem[14307] <= 16'hFFFF;
rommem[14308] <= 16'hFFFF;
rommem[14309] <= 16'hFFFF;
rommem[14310] <= 16'hFFFF;
rommem[14311] <= 16'hFFFF;
rommem[14312] <= 16'hFFFF;
rommem[14313] <= 16'hFFFF;
rommem[14314] <= 16'hFFFF;
rommem[14315] <= 16'hFFFF;
rommem[14316] <= 16'hFFFF;
rommem[14317] <= 16'hFFFF;
rommem[14318] <= 16'hFFFF;
rommem[14319] <= 16'hFFFF;
rommem[14320] <= 16'hFFFF;
rommem[14321] <= 16'hFFFF;
rommem[14322] <= 16'hFFFF;
rommem[14323] <= 16'hFFFF;
rommem[14324] <= 16'hFFFF;
rommem[14325] <= 16'hFFFF;
rommem[14326] <= 16'hFFFF;
rommem[14327] <= 16'hFFFF;
rommem[14328] <= 16'hFFFF;
rommem[14329] <= 16'hFFFF;
rommem[14330] <= 16'hFFFF;
rommem[14331] <= 16'hFFFF;
rommem[14332] <= 16'hFFFF;
rommem[14333] <= 16'hFFFF;
rommem[14334] <= 16'hFFFF;
rommem[14335] <= 16'hFFFF;
rommem[14336] <= 16'hFFFF;
rommem[14337] <= 16'hFFFF;
rommem[14338] <= 16'hFFFF;
rommem[14339] <= 16'hFFFF;
rommem[14340] <= 16'hFFFF;
rommem[14341] <= 16'hFFFF;
rommem[14342] <= 16'hFFFF;
rommem[14343] <= 16'hFFFF;
rommem[14344] <= 16'hFFFF;
rommem[14345] <= 16'hFFFF;
rommem[14346] <= 16'hFFFF;
rommem[14347] <= 16'hFFFF;
rommem[14348] <= 16'hFFFF;
rommem[14349] <= 16'hFFFF;
rommem[14350] <= 16'hFFFF;
rommem[14351] <= 16'hFFFF;
rommem[14352] <= 16'hFFFF;
rommem[14353] <= 16'hFFFF;
rommem[14354] <= 16'hFFFF;
rommem[14355] <= 16'hFFFF;
rommem[14356] <= 16'hFFFF;
rommem[14357] <= 16'hFFFF;
rommem[14358] <= 16'hFFFF;
rommem[14359] <= 16'hFFFF;
rommem[14360] <= 16'hFFFF;
rommem[14361] <= 16'hFFFF;
rommem[14362] <= 16'hFFFF;
rommem[14363] <= 16'hFFFF;
rommem[14364] <= 16'hFFFF;
rommem[14365] <= 16'hFFFF;
rommem[14366] <= 16'hFFFF;
rommem[14367] <= 16'hFFFF;
rommem[14368] <= 16'hFFFF;
rommem[14369] <= 16'hFFFF;
rommem[14370] <= 16'hFFFF;
rommem[14371] <= 16'hFFFF;
rommem[14372] <= 16'hFFFF;
rommem[14373] <= 16'hFFFF;
rommem[14374] <= 16'hFFFF;
rommem[14375] <= 16'hFFFF;
rommem[14376] <= 16'hFFFF;
rommem[14377] <= 16'hFFFF;
rommem[14378] <= 16'hFFFF;
rommem[14379] <= 16'hFFFF;
rommem[14380] <= 16'hFFFF;
rommem[14381] <= 16'hFFFF;
rommem[14382] <= 16'hFFFF;
rommem[14383] <= 16'hFFFF;
rommem[14384] <= 16'hFFFF;
rommem[14385] <= 16'hFFFF;
rommem[14386] <= 16'hFFFF;
rommem[14387] <= 16'hFFFF;
rommem[14388] <= 16'hFFFF;
rommem[14389] <= 16'hFFFF;
rommem[14390] <= 16'hFFFF;
rommem[14391] <= 16'hFFFF;
rommem[14392] <= 16'hFFFF;
rommem[14393] <= 16'hFFFF;
rommem[14394] <= 16'hFFFF;
rommem[14395] <= 16'hFFFF;
rommem[14396] <= 16'hFFFF;
rommem[14397] <= 16'hFFFF;
rommem[14398] <= 16'hFFFF;
rommem[14399] <= 16'hFFFF;
rommem[14400] <= 16'hFFFF;
rommem[14401] <= 16'hFFFF;
rommem[14402] <= 16'hFFFF;
rommem[14403] <= 16'hFFFF;
rommem[14404] <= 16'hFFFF;
rommem[14405] <= 16'hFFFF;
rommem[14406] <= 16'hFFFF;
rommem[14407] <= 16'hFFFF;
rommem[14408] <= 16'hFFFF;
rommem[14409] <= 16'hFFFF;
rommem[14410] <= 16'hFFFF;
rommem[14411] <= 16'hFFFF;
rommem[14412] <= 16'hFFFF;
rommem[14413] <= 16'hFFFF;
rommem[14414] <= 16'hFFFF;
rommem[14415] <= 16'hFFFF;
rommem[14416] <= 16'hFFFF;
rommem[14417] <= 16'hFFFF;
rommem[14418] <= 16'hFFFF;
rommem[14419] <= 16'hFFFF;
rommem[14420] <= 16'hFFFF;
rommem[14421] <= 16'hFFFF;
rommem[14422] <= 16'hFFFF;
rommem[14423] <= 16'hFFFF;
rommem[14424] <= 16'hFFFF;
rommem[14425] <= 16'hFFFF;
rommem[14426] <= 16'hFFFF;
rommem[14427] <= 16'hFFFF;
rommem[14428] <= 16'hFFFF;
rommem[14429] <= 16'hFFFF;
rommem[14430] <= 16'hFFFF;
rommem[14431] <= 16'hFFFF;
rommem[14432] <= 16'hFFFF;
rommem[14433] <= 16'hFFFF;
rommem[14434] <= 16'hFFFF;
rommem[14435] <= 16'hFFFF;
rommem[14436] <= 16'hFFFF;
rommem[14437] <= 16'hFFFF;
rommem[14438] <= 16'hFFFF;
rommem[14439] <= 16'hFFFF;
rommem[14440] <= 16'hFFFF;
rommem[14441] <= 16'hFFFF;
rommem[14442] <= 16'hFFFF;
rommem[14443] <= 16'hFFFF;
rommem[14444] <= 16'hFFFF;
rommem[14445] <= 16'hFFFF;
rommem[14446] <= 16'hFFFF;
rommem[14447] <= 16'hFFFF;
rommem[14448] <= 16'hFFFF;
rommem[14449] <= 16'hFFFF;
rommem[14450] <= 16'hFFFF;
rommem[14451] <= 16'hFFFF;
rommem[14452] <= 16'hFFFF;
rommem[14453] <= 16'hFFFF;
rommem[14454] <= 16'hFFFF;
rommem[14455] <= 16'hFFFF;
rommem[14456] <= 16'hFFFF;
rommem[14457] <= 16'hFFFF;
rommem[14458] <= 16'hFFFF;
rommem[14459] <= 16'hFFFF;
rommem[14460] <= 16'hFFFF;
rommem[14461] <= 16'hFFFF;
rommem[14462] <= 16'hFFFF;
rommem[14463] <= 16'hFFFF;
rommem[14464] <= 16'hFFFF;
rommem[14465] <= 16'hFFFF;
rommem[14466] <= 16'hFFFF;
rommem[14467] <= 16'hFFFF;
rommem[14468] <= 16'hFFFF;
rommem[14469] <= 16'hFFFF;
rommem[14470] <= 16'hFFFF;
rommem[14471] <= 16'hFFFF;
rommem[14472] <= 16'hFFFF;
rommem[14473] <= 16'hFFFF;
rommem[14474] <= 16'hFFFF;
rommem[14475] <= 16'hFFFF;
rommem[14476] <= 16'hFFFF;
rommem[14477] <= 16'hFFFF;
rommem[14478] <= 16'hFFFF;
rommem[14479] <= 16'hFFFF;
rommem[14480] <= 16'hFFFF;
rommem[14481] <= 16'hFFFF;
rommem[14482] <= 16'hFFFF;
rommem[14483] <= 16'hFFFF;
rommem[14484] <= 16'hFFFF;
rommem[14485] <= 16'hFFFF;
rommem[14486] <= 16'hFFFF;
rommem[14487] <= 16'hFFFF;
rommem[14488] <= 16'hFFFF;
rommem[14489] <= 16'hFFFF;
rommem[14490] <= 16'hFFFF;
rommem[14491] <= 16'hFFFF;
rommem[14492] <= 16'hFFFF;
rommem[14493] <= 16'hFFFF;
rommem[14494] <= 16'hFFFF;
rommem[14495] <= 16'hFFFF;
rommem[14496] <= 16'hFFFF;
rommem[14497] <= 16'hFFFF;
rommem[14498] <= 16'hFFFF;
rommem[14499] <= 16'hFFFF;
rommem[14500] <= 16'hFFFF;
rommem[14501] <= 16'hFFFF;
rommem[14502] <= 16'hFFFF;
rommem[14503] <= 16'hFFFF;
rommem[14504] <= 16'hFFFF;
rommem[14505] <= 16'hFFFF;
rommem[14506] <= 16'hFFFF;
rommem[14507] <= 16'hFFFF;
rommem[14508] <= 16'hFFFF;
rommem[14509] <= 16'hFFFF;
rommem[14510] <= 16'hFFFF;
rommem[14511] <= 16'hFFFF;
rommem[14512] <= 16'hFFFF;
rommem[14513] <= 16'hFFFF;
rommem[14514] <= 16'hFFFF;
rommem[14515] <= 16'hFFFF;
rommem[14516] <= 16'hFFFF;
rommem[14517] <= 16'hFFFF;
rommem[14518] <= 16'hFFFF;
rommem[14519] <= 16'hFFFF;
rommem[14520] <= 16'hFFFF;
rommem[14521] <= 16'hFFFF;
rommem[14522] <= 16'hFFFF;
rommem[14523] <= 16'hFFFF;
rommem[14524] <= 16'hFFFF;
rommem[14525] <= 16'hFFFF;
rommem[14526] <= 16'hFFFF;
rommem[14527] <= 16'hFFFF;
rommem[14528] <= 16'hFFFF;
rommem[14529] <= 16'hFFFF;
rommem[14530] <= 16'hFFFF;
rommem[14531] <= 16'hFFFF;
rommem[14532] <= 16'hFFFF;
rommem[14533] <= 16'hFFFF;
rommem[14534] <= 16'hFFFF;
rommem[14535] <= 16'hFFFF;
rommem[14536] <= 16'hFFFF;
rommem[14537] <= 16'hFFFF;
rommem[14538] <= 16'hFFFF;
rommem[14539] <= 16'hFFFF;
rommem[14540] <= 16'hFFFF;
rommem[14541] <= 16'hFFFF;
rommem[14542] <= 16'hFFFF;
rommem[14543] <= 16'hFFFF;
rommem[14544] <= 16'hFFFF;
rommem[14545] <= 16'hFFFF;
rommem[14546] <= 16'hFFFF;
rommem[14547] <= 16'hFFFF;
rommem[14548] <= 16'hFFFF;
rommem[14549] <= 16'hFFFF;
rommem[14550] <= 16'hFFFF;
rommem[14551] <= 16'hFFFF;
rommem[14552] <= 16'hFFFF;
rommem[14553] <= 16'hFFFF;
rommem[14554] <= 16'hFFFF;
rommem[14555] <= 16'hFFFF;
rommem[14556] <= 16'hFFFF;
rommem[14557] <= 16'hFFFF;
rommem[14558] <= 16'hFFFF;
rommem[14559] <= 16'hFFFF;
rommem[14560] <= 16'hFFFF;
rommem[14561] <= 16'hFFFF;
rommem[14562] <= 16'hFFFF;
rommem[14563] <= 16'hFFFF;
rommem[14564] <= 16'hFFFF;
rommem[14565] <= 16'hFFFF;
rommem[14566] <= 16'hFFFF;
rommem[14567] <= 16'hFFFF;
rommem[14568] <= 16'hFFFF;
rommem[14569] <= 16'hFFFF;
rommem[14570] <= 16'hFFFF;
rommem[14571] <= 16'hFFFF;
rommem[14572] <= 16'hFFFF;
rommem[14573] <= 16'hFFFF;
rommem[14574] <= 16'hFFFF;
rommem[14575] <= 16'hFFFF;
rommem[14576] <= 16'hFFFF;
rommem[14577] <= 16'hFFFF;
rommem[14578] <= 16'hFFFF;
rommem[14579] <= 16'hFFFF;
rommem[14580] <= 16'hFFFF;
rommem[14581] <= 16'hFFFF;
rommem[14582] <= 16'hFFFF;
rommem[14583] <= 16'hFFFF;
rommem[14584] <= 16'hFFFF;
rommem[14585] <= 16'hFFFF;
rommem[14586] <= 16'hFFFF;
rommem[14587] <= 16'hFFFF;
rommem[14588] <= 16'hFFFF;
rommem[14589] <= 16'hFFFF;
rommem[14590] <= 16'hFFFF;
rommem[14591] <= 16'hFFFF;
rommem[14592] <= 16'hFFFF;
rommem[14593] <= 16'hFFFF;
rommem[14594] <= 16'hFFFF;
rommem[14595] <= 16'hFFFF;
rommem[14596] <= 16'hFFFF;
rommem[14597] <= 16'hFFFF;
rommem[14598] <= 16'hFFFF;
rommem[14599] <= 16'hFFFF;
rommem[14600] <= 16'hFFFF;
rommem[14601] <= 16'hFFFF;
rommem[14602] <= 16'hFFFF;
rommem[14603] <= 16'hFFFF;
rommem[14604] <= 16'hFFFF;
rommem[14605] <= 16'hFFFF;
rommem[14606] <= 16'hFFFF;
rommem[14607] <= 16'hFFFF;
rommem[14608] <= 16'hFFFF;
rommem[14609] <= 16'hFFFF;
rommem[14610] <= 16'hFFFF;
rommem[14611] <= 16'hFFFF;
rommem[14612] <= 16'hFFFF;
rommem[14613] <= 16'hFFFF;
rommem[14614] <= 16'hFFFF;
rommem[14615] <= 16'hFFFF;
rommem[14616] <= 16'hFFFF;
rommem[14617] <= 16'hFFFF;
rommem[14618] <= 16'hFFFF;
rommem[14619] <= 16'hFFFF;
rommem[14620] <= 16'hFFFF;
rommem[14621] <= 16'hFFFF;
rommem[14622] <= 16'hFFFF;
rommem[14623] <= 16'hFFFF;
rommem[14624] <= 16'hFFFF;
rommem[14625] <= 16'hFFFF;
rommem[14626] <= 16'hFFFF;
rommem[14627] <= 16'hFFFF;
rommem[14628] <= 16'hFFFF;
rommem[14629] <= 16'hFFFF;
rommem[14630] <= 16'hFFFF;
rommem[14631] <= 16'hFFFF;
rommem[14632] <= 16'hFFFF;
rommem[14633] <= 16'hFFFF;
rommem[14634] <= 16'hFFFF;
rommem[14635] <= 16'hFFFF;
rommem[14636] <= 16'hFFFF;
rommem[14637] <= 16'hFFFF;
rommem[14638] <= 16'hFFFF;
rommem[14639] <= 16'hFFFF;
rommem[14640] <= 16'hFFFF;
rommem[14641] <= 16'hFFFF;
rommem[14642] <= 16'hFFFF;
rommem[14643] <= 16'hFFFF;
rommem[14644] <= 16'hFFFF;
rommem[14645] <= 16'hFFFF;
rommem[14646] <= 16'hFFFF;
rommem[14647] <= 16'hFFFF;
rommem[14648] <= 16'hFFFF;
rommem[14649] <= 16'hFFFF;
rommem[14650] <= 16'hFFFF;
rommem[14651] <= 16'hFFFF;
rommem[14652] <= 16'hFFFF;
rommem[14653] <= 16'hFFFF;
rommem[14654] <= 16'hFFFF;
rommem[14655] <= 16'hFFFF;
rommem[14656] <= 16'hFFFF;
rommem[14657] <= 16'hFFFF;
rommem[14658] <= 16'hFFFF;
rommem[14659] <= 16'hFFFF;
rommem[14660] <= 16'hFFFF;
rommem[14661] <= 16'hFFFF;
rommem[14662] <= 16'hFFFF;
rommem[14663] <= 16'hFFFF;
rommem[14664] <= 16'hFFFF;
rommem[14665] <= 16'hFFFF;
rommem[14666] <= 16'hFFFF;
rommem[14667] <= 16'hFFFF;
rommem[14668] <= 16'hFFFF;
rommem[14669] <= 16'hFFFF;
rommem[14670] <= 16'hFFFF;
rommem[14671] <= 16'hFFFF;
rommem[14672] <= 16'hFFFF;
rommem[14673] <= 16'hFFFF;
rommem[14674] <= 16'hFFFF;
rommem[14675] <= 16'hFFFF;
rommem[14676] <= 16'hFFFF;
rommem[14677] <= 16'hFFFF;
rommem[14678] <= 16'hFFFF;
rommem[14679] <= 16'hFFFF;
rommem[14680] <= 16'hFFFF;
rommem[14681] <= 16'hFFFF;
rommem[14682] <= 16'hFFFF;
rommem[14683] <= 16'hFFFF;
rommem[14684] <= 16'hFFFF;
rommem[14685] <= 16'hFFFF;
rommem[14686] <= 16'hFFFF;
rommem[14687] <= 16'hFFFF;
rommem[14688] <= 16'hFFFF;
rommem[14689] <= 16'hFFFF;
rommem[14690] <= 16'hFFFF;
rommem[14691] <= 16'hFFFF;
rommem[14692] <= 16'hFFFF;
rommem[14693] <= 16'hFFFF;
rommem[14694] <= 16'hFFFF;
rommem[14695] <= 16'hFFFF;
rommem[14696] <= 16'hFFFF;
rommem[14697] <= 16'hFFFF;
rommem[14698] <= 16'hFFFF;
rommem[14699] <= 16'hFFFF;
rommem[14700] <= 16'hFFFF;
rommem[14701] <= 16'hFFFF;
rommem[14702] <= 16'hFFFF;
rommem[14703] <= 16'hFFFF;
rommem[14704] <= 16'hFFFF;
rommem[14705] <= 16'hFFFF;
rommem[14706] <= 16'hFFFF;
rommem[14707] <= 16'hFFFF;
rommem[14708] <= 16'hFFFF;
rommem[14709] <= 16'hFFFF;
rommem[14710] <= 16'hFFFF;
rommem[14711] <= 16'hFFFF;
rommem[14712] <= 16'hFFFF;
rommem[14713] <= 16'hFFFF;
rommem[14714] <= 16'hFFFF;
rommem[14715] <= 16'hFFFF;
rommem[14716] <= 16'hFFFF;
rommem[14717] <= 16'hFFFF;
rommem[14718] <= 16'hFFFF;
rommem[14719] <= 16'hFFFF;
rommem[14720] <= 16'hFFFF;
rommem[14721] <= 16'hFFFF;
rommem[14722] <= 16'hFFFF;
rommem[14723] <= 16'hFFFF;
rommem[14724] <= 16'hFFFF;
rommem[14725] <= 16'hFFFF;
rommem[14726] <= 16'hFFFF;
rommem[14727] <= 16'hFFFF;
rommem[14728] <= 16'hFFFF;
rommem[14729] <= 16'hFFFF;
rommem[14730] <= 16'hFFFF;
rommem[14731] <= 16'hFFFF;
rommem[14732] <= 16'hFFFF;
rommem[14733] <= 16'hFFFF;
rommem[14734] <= 16'hFFFF;
rommem[14735] <= 16'hFFFF;
rommem[14736] <= 16'hFFFF;
rommem[14737] <= 16'hFFFF;
rommem[14738] <= 16'hFFFF;
rommem[14739] <= 16'hFFFF;
rommem[14740] <= 16'hFFFF;
rommem[14741] <= 16'hFFFF;
rommem[14742] <= 16'hFFFF;
rommem[14743] <= 16'hFFFF;
rommem[14744] <= 16'hFFFF;
rommem[14745] <= 16'hFFFF;
rommem[14746] <= 16'hFFFF;
rommem[14747] <= 16'hFFFF;
rommem[14748] <= 16'hFFFF;
rommem[14749] <= 16'hFFFF;
rommem[14750] <= 16'hFFFF;
rommem[14751] <= 16'hFFFF;
rommem[14752] <= 16'hFFFF;
rommem[14753] <= 16'hFFFF;
rommem[14754] <= 16'hFFFF;
rommem[14755] <= 16'hFFFF;
rommem[14756] <= 16'hFFFF;
rommem[14757] <= 16'hFFFF;
rommem[14758] <= 16'hFFFF;
rommem[14759] <= 16'hFFFF;
rommem[14760] <= 16'hFFFF;
rommem[14761] <= 16'hFFFF;
rommem[14762] <= 16'hFFFF;
rommem[14763] <= 16'hFFFF;
rommem[14764] <= 16'hFFFF;
rommem[14765] <= 16'hFFFF;
rommem[14766] <= 16'hFFFF;
rommem[14767] <= 16'hFFFF;
rommem[14768] <= 16'hFFFF;
rommem[14769] <= 16'hFFFF;
rommem[14770] <= 16'hFFFF;
rommem[14771] <= 16'hFFFF;
rommem[14772] <= 16'hFFFF;
rommem[14773] <= 16'hFFFF;
rommem[14774] <= 16'hFFFF;
rommem[14775] <= 16'hFFFF;
rommem[14776] <= 16'hFFFF;
rommem[14777] <= 16'hFFFF;
rommem[14778] <= 16'hFFFF;
rommem[14779] <= 16'hFFFF;
rommem[14780] <= 16'hFFFF;
rommem[14781] <= 16'hFFFF;
rommem[14782] <= 16'hFFFF;
rommem[14783] <= 16'hFFFF;
rommem[14784] <= 16'hFFFF;
rommem[14785] <= 16'hFFFF;
rommem[14786] <= 16'hFFFF;
rommem[14787] <= 16'hFFFF;
rommem[14788] <= 16'hFFFF;
rommem[14789] <= 16'hFFFF;
rommem[14790] <= 16'hFFFF;
rommem[14791] <= 16'hFFFF;
rommem[14792] <= 16'hFFFF;
rommem[14793] <= 16'hFFFF;
rommem[14794] <= 16'hFFFF;
rommem[14795] <= 16'hFFFF;
rommem[14796] <= 16'hFFFF;
rommem[14797] <= 16'hFFFF;
rommem[14798] <= 16'hFFFF;
rommem[14799] <= 16'hFFFF;
rommem[14800] <= 16'hFFFF;
rommem[14801] <= 16'hFFFF;
rommem[14802] <= 16'hFFFF;
rommem[14803] <= 16'hFFFF;
rommem[14804] <= 16'hFFFF;
rommem[14805] <= 16'hFFFF;
rommem[14806] <= 16'hFFFF;
rommem[14807] <= 16'hFFFF;
rommem[14808] <= 16'hFFFF;
rommem[14809] <= 16'hFFFF;
rommem[14810] <= 16'hFFFF;
rommem[14811] <= 16'hFFFF;
rommem[14812] <= 16'hFFFF;
rommem[14813] <= 16'hFFFF;
rommem[14814] <= 16'hFFFF;
rommem[14815] <= 16'hFFFF;
rommem[14816] <= 16'hFFFF;
rommem[14817] <= 16'hFFFF;
rommem[14818] <= 16'hFFFF;
rommem[14819] <= 16'hFFFF;
rommem[14820] <= 16'hFFFF;
rommem[14821] <= 16'hFFFF;
rommem[14822] <= 16'hFFFF;
rommem[14823] <= 16'hFFFF;
rommem[14824] <= 16'hFFFF;
rommem[14825] <= 16'hFFFF;
rommem[14826] <= 16'hFFFF;
rommem[14827] <= 16'hFFFF;
rommem[14828] <= 16'hFFFF;
rommem[14829] <= 16'hFFFF;
rommem[14830] <= 16'hFFFF;
rommem[14831] <= 16'hFFFF;
rommem[14832] <= 16'hFFFF;
rommem[14833] <= 16'hFFFF;
rommem[14834] <= 16'hFFFF;
rommem[14835] <= 16'hFFFF;
rommem[14836] <= 16'hFFFF;
rommem[14837] <= 16'hFFFF;
rommem[14838] <= 16'hFFFF;
rommem[14839] <= 16'hFFFF;
rommem[14840] <= 16'hFFFF;
rommem[14841] <= 16'hFFFF;
rommem[14842] <= 16'hFFFF;
rommem[14843] <= 16'hFFFF;
rommem[14844] <= 16'hFFFF;
rommem[14845] <= 16'hFFFF;
rommem[14846] <= 16'hFFFF;
rommem[14847] <= 16'hFFFF;
rommem[14848] <= 16'hFFFF;
rommem[14849] <= 16'hFFFF;
rommem[14850] <= 16'hFFFF;
rommem[14851] <= 16'hFFFF;
rommem[14852] <= 16'hFFFF;
rommem[14853] <= 16'hFFFF;
rommem[14854] <= 16'hFFFF;
rommem[14855] <= 16'hFFFF;
rommem[14856] <= 16'hFFFF;
rommem[14857] <= 16'hFFFF;
rommem[14858] <= 16'hFFFF;
rommem[14859] <= 16'hFFFF;
rommem[14860] <= 16'hFFFF;
rommem[14861] <= 16'hFFFF;
rommem[14862] <= 16'hFFFF;
rommem[14863] <= 16'hFFFF;
rommem[14864] <= 16'hFFFF;
rommem[14865] <= 16'hFFFF;
rommem[14866] <= 16'hFFFF;
rommem[14867] <= 16'hFFFF;
rommem[14868] <= 16'hFFFF;
rommem[14869] <= 16'hFFFF;
rommem[14870] <= 16'hFFFF;
rommem[14871] <= 16'hFFFF;
rommem[14872] <= 16'hFFFF;
rommem[14873] <= 16'hFFFF;
rommem[14874] <= 16'hFFFF;
rommem[14875] <= 16'hFFFF;
rommem[14876] <= 16'hFFFF;
rommem[14877] <= 16'hFFFF;
rommem[14878] <= 16'hFFFF;
rommem[14879] <= 16'hFFFF;
rommem[14880] <= 16'hFFFF;
rommem[14881] <= 16'hFFFF;
rommem[14882] <= 16'hFFFF;
rommem[14883] <= 16'hFFFF;
rommem[14884] <= 16'hFFFF;
rommem[14885] <= 16'hFFFF;
rommem[14886] <= 16'hFFFF;
rommem[14887] <= 16'hFFFF;
rommem[14888] <= 16'hFFFF;
rommem[14889] <= 16'hFFFF;
rommem[14890] <= 16'hFFFF;
rommem[14891] <= 16'hFFFF;
rommem[14892] <= 16'hFFFF;
rommem[14893] <= 16'hFFFF;
rommem[14894] <= 16'hFFFF;
rommem[14895] <= 16'hFFFF;
rommem[14896] <= 16'hFFFF;
rommem[14897] <= 16'hFFFF;
rommem[14898] <= 16'hFFFF;
rommem[14899] <= 16'hFFFF;
rommem[14900] <= 16'hFFFF;
rommem[14901] <= 16'hFFFF;
rommem[14902] <= 16'hFFFF;
rommem[14903] <= 16'hFFFF;
rommem[14904] <= 16'hFFFF;
rommem[14905] <= 16'hFFFF;
rommem[14906] <= 16'hFFFF;
rommem[14907] <= 16'hFFFF;
rommem[14908] <= 16'hFFFF;
rommem[14909] <= 16'hFFFF;
rommem[14910] <= 16'hFFFF;
rommem[14911] <= 16'hFFFF;
rommem[14912] <= 16'hFFFF;
rommem[14913] <= 16'hFFFF;
rommem[14914] <= 16'hFFFF;
rommem[14915] <= 16'hFFFF;
rommem[14916] <= 16'hFFFF;
rommem[14917] <= 16'hFFFF;
rommem[14918] <= 16'hFFFF;
rommem[14919] <= 16'hFFFF;
rommem[14920] <= 16'hFFFF;
rommem[14921] <= 16'hFFFF;
rommem[14922] <= 16'hFFFF;
rommem[14923] <= 16'hFFFF;
rommem[14924] <= 16'hFFFF;
rommem[14925] <= 16'hFFFF;
rommem[14926] <= 16'hFFFF;
rommem[14927] <= 16'hFFFF;
rommem[14928] <= 16'hFFFF;
rommem[14929] <= 16'hFFFF;
rommem[14930] <= 16'hFFFF;
rommem[14931] <= 16'hFFFF;
rommem[14932] <= 16'hFFFF;
rommem[14933] <= 16'hFFFF;
rommem[14934] <= 16'hFFFF;
rommem[14935] <= 16'hFFFF;
rommem[14936] <= 16'hFFFF;
rommem[14937] <= 16'hFFFF;
rommem[14938] <= 16'hFFFF;
rommem[14939] <= 16'hFFFF;
rommem[14940] <= 16'hFFFF;
rommem[14941] <= 16'hFFFF;
rommem[14942] <= 16'hFFFF;
rommem[14943] <= 16'hFFFF;
rommem[14944] <= 16'hFFFF;
rommem[14945] <= 16'hFFFF;
rommem[14946] <= 16'hFFFF;
rommem[14947] <= 16'hFFFF;
rommem[14948] <= 16'hFFFF;
rommem[14949] <= 16'hFFFF;
rommem[14950] <= 16'hFFFF;
rommem[14951] <= 16'hFFFF;
rommem[14952] <= 16'hFFFF;
rommem[14953] <= 16'hFFFF;
rommem[14954] <= 16'hFFFF;
rommem[14955] <= 16'hFFFF;
rommem[14956] <= 16'hFFFF;
rommem[14957] <= 16'hFFFF;
rommem[14958] <= 16'hFFFF;
rommem[14959] <= 16'hFFFF;
rommem[14960] <= 16'hFFFF;
rommem[14961] <= 16'hFFFF;
rommem[14962] <= 16'hFFFF;
rommem[14963] <= 16'hFFFF;
rommem[14964] <= 16'hFFFF;
rommem[14965] <= 16'hFFFF;
rommem[14966] <= 16'hFFFF;
rommem[14967] <= 16'hFFFF;
rommem[14968] <= 16'hFFFF;
rommem[14969] <= 16'hFFFF;
rommem[14970] <= 16'hFFFF;
rommem[14971] <= 16'hFFFF;
rommem[14972] <= 16'hFFFF;
rommem[14973] <= 16'hFFFF;
rommem[14974] <= 16'hFFFF;
rommem[14975] <= 16'hFFFF;
rommem[14976] <= 16'hFFFF;
rommem[14977] <= 16'hFFFF;
rommem[14978] <= 16'hFFFF;
rommem[14979] <= 16'hFFFF;
rommem[14980] <= 16'hFFFF;
rommem[14981] <= 16'hFFFF;
rommem[14982] <= 16'hFFFF;
rommem[14983] <= 16'hFFFF;
rommem[14984] <= 16'hFFFF;
rommem[14985] <= 16'hFFFF;
rommem[14986] <= 16'hFFFF;
rommem[14987] <= 16'hFFFF;
rommem[14988] <= 16'hFFFF;
rommem[14989] <= 16'hFFFF;
rommem[14990] <= 16'hFFFF;
rommem[14991] <= 16'hFFFF;
rommem[14992] <= 16'hFFFF;
rommem[14993] <= 16'hFFFF;
rommem[14994] <= 16'hFFFF;
rommem[14995] <= 16'hFFFF;
rommem[14996] <= 16'hFFFF;
rommem[14997] <= 16'hFFFF;
rommem[14998] <= 16'hFFFF;
rommem[14999] <= 16'hFFFF;
rommem[15000] <= 16'hFFFF;
rommem[15001] <= 16'hFFFF;
rommem[15002] <= 16'hFFFF;
rommem[15003] <= 16'hFFFF;
rommem[15004] <= 16'hFFFF;
rommem[15005] <= 16'hFFFF;
rommem[15006] <= 16'hFFFF;
rommem[15007] <= 16'hFFFF;
rommem[15008] <= 16'hFFFF;
rommem[15009] <= 16'hFFFF;
rommem[15010] <= 16'hFFFF;
rommem[15011] <= 16'hFFFF;
rommem[15012] <= 16'hFFFF;
rommem[15013] <= 16'hFFFF;
rommem[15014] <= 16'hFFFF;
rommem[15015] <= 16'hFFFF;
rommem[15016] <= 16'hFFFF;
rommem[15017] <= 16'hFFFF;
rommem[15018] <= 16'hFFFF;
rommem[15019] <= 16'hFFFF;
rommem[15020] <= 16'hFFFF;
rommem[15021] <= 16'hFFFF;
rommem[15022] <= 16'hFFFF;
rommem[15023] <= 16'hFFFF;
rommem[15024] <= 16'hFFFF;
rommem[15025] <= 16'hFFFF;
rommem[15026] <= 16'hFFFF;
rommem[15027] <= 16'hFFFF;
rommem[15028] <= 16'hFFFF;
rommem[15029] <= 16'hFFFF;
rommem[15030] <= 16'hFFFF;
rommem[15031] <= 16'hFFFF;
rommem[15032] <= 16'hFFFF;
rommem[15033] <= 16'hFFFF;
rommem[15034] <= 16'hFFFF;
rommem[15035] <= 16'hFFFF;
rommem[15036] <= 16'hFFFF;
rommem[15037] <= 16'hFFFF;
rommem[15038] <= 16'hFFFF;
rommem[15039] <= 16'hFFFF;
rommem[15040] <= 16'hFFFF;
rommem[15041] <= 16'hFFFF;
rommem[15042] <= 16'hFFFF;
rommem[15043] <= 16'hFFFF;
rommem[15044] <= 16'hFFFF;
rommem[15045] <= 16'hFFFF;
rommem[15046] <= 16'hFFFF;
rommem[15047] <= 16'hFFFF;
rommem[15048] <= 16'hFFFF;
rommem[15049] <= 16'hFFFF;
rommem[15050] <= 16'hFFFF;
rommem[15051] <= 16'hFFFF;
rommem[15052] <= 16'hFFFF;
rommem[15053] <= 16'hFFFF;
rommem[15054] <= 16'hFFFF;
rommem[15055] <= 16'hFFFF;
rommem[15056] <= 16'hFFFF;
rommem[15057] <= 16'hFFFF;
rommem[15058] <= 16'hFFFF;
rommem[15059] <= 16'hFFFF;
rommem[15060] <= 16'hFFFF;
rommem[15061] <= 16'hFFFF;
rommem[15062] <= 16'hFFFF;
rommem[15063] <= 16'hFFFF;
rommem[15064] <= 16'hFFFF;
rommem[15065] <= 16'hFFFF;
rommem[15066] <= 16'hFFFF;
rommem[15067] <= 16'hFFFF;
rommem[15068] <= 16'hFFFF;
rommem[15069] <= 16'hFFFF;
rommem[15070] <= 16'hFFFF;
rommem[15071] <= 16'hFFFF;
rommem[15072] <= 16'hFFFF;
rommem[15073] <= 16'hFFFF;
rommem[15074] <= 16'hFFFF;
rommem[15075] <= 16'hFFFF;
rommem[15076] <= 16'hFFFF;
rommem[15077] <= 16'hFFFF;
rommem[15078] <= 16'hFFFF;
rommem[15079] <= 16'hFFFF;
rommem[15080] <= 16'hFFFF;
rommem[15081] <= 16'hFFFF;
rommem[15082] <= 16'hFFFF;
rommem[15083] <= 16'hFFFF;
rommem[15084] <= 16'hFFFF;
rommem[15085] <= 16'hFFFF;
rommem[15086] <= 16'hFFFF;
rommem[15087] <= 16'hFFFF;
rommem[15088] <= 16'hFFFF;
rommem[15089] <= 16'hFFFF;
rommem[15090] <= 16'hFFFF;
rommem[15091] <= 16'hFFFF;
rommem[15092] <= 16'hFFFF;
rommem[15093] <= 16'hFFFF;
rommem[15094] <= 16'hFFFF;
rommem[15095] <= 16'hFFFF;
rommem[15096] <= 16'hFFFF;
rommem[15097] <= 16'hFFFF;
rommem[15098] <= 16'hFFFF;
rommem[15099] <= 16'hFFFF;
rommem[15100] <= 16'hFFFF;
rommem[15101] <= 16'hFFFF;
rommem[15102] <= 16'hFFFF;
rommem[15103] <= 16'hFFFF;
rommem[15104] <= 16'hFFFF;
rommem[15105] <= 16'hFFFF;
rommem[15106] <= 16'hFFFF;
rommem[15107] <= 16'hFFFF;
rommem[15108] <= 16'hFFFF;
rommem[15109] <= 16'hFFFF;
rommem[15110] <= 16'hFFFF;
rommem[15111] <= 16'hFFFF;
rommem[15112] <= 16'hFFFF;
rommem[15113] <= 16'hFFFF;
rommem[15114] <= 16'hFFFF;
rommem[15115] <= 16'hFFFF;
rommem[15116] <= 16'hFFFF;
rommem[15117] <= 16'hFFFF;
rommem[15118] <= 16'hFFFF;
rommem[15119] <= 16'hFFFF;
rommem[15120] <= 16'hFFFF;
rommem[15121] <= 16'hFFFF;
rommem[15122] <= 16'hFFFF;
rommem[15123] <= 16'hFFFF;
rommem[15124] <= 16'hFFFF;
rommem[15125] <= 16'hFFFF;
rommem[15126] <= 16'hFFFF;
rommem[15127] <= 16'hFFFF;
rommem[15128] <= 16'hFFFF;
rommem[15129] <= 16'hFFFF;
rommem[15130] <= 16'hFFFF;
rommem[15131] <= 16'hFFFF;
rommem[15132] <= 16'hFFFF;
rommem[15133] <= 16'hFFFF;
rommem[15134] <= 16'hFFFF;
rommem[15135] <= 16'hFFFF;
rommem[15136] <= 16'hFFFF;
rommem[15137] <= 16'hFFFF;
rommem[15138] <= 16'hFFFF;
rommem[15139] <= 16'hFFFF;
rommem[15140] <= 16'hFFFF;
rommem[15141] <= 16'hFFFF;
rommem[15142] <= 16'hFFFF;
rommem[15143] <= 16'hFFFF;
rommem[15144] <= 16'hFFFF;
rommem[15145] <= 16'hFFFF;
rommem[15146] <= 16'hFFFF;
rommem[15147] <= 16'hFFFF;
rommem[15148] <= 16'hFFFF;
rommem[15149] <= 16'hFFFF;
rommem[15150] <= 16'hFFFF;
rommem[15151] <= 16'hFFFF;
rommem[15152] <= 16'hFFFF;
rommem[15153] <= 16'hFFFF;
rommem[15154] <= 16'hFFFF;
rommem[15155] <= 16'hFFFF;
rommem[15156] <= 16'hFFFF;
rommem[15157] <= 16'hFFFF;
rommem[15158] <= 16'hFFFF;
rommem[15159] <= 16'hFFFF;
rommem[15160] <= 16'hFFFF;
rommem[15161] <= 16'hFFFF;
rommem[15162] <= 16'hFFFF;
rommem[15163] <= 16'hFFFF;
rommem[15164] <= 16'hFFFF;
rommem[15165] <= 16'hFFFF;
rommem[15166] <= 16'hFFFF;
rommem[15167] <= 16'hFFFF;
rommem[15168] <= 16'hFFFF;
rommem[15169] <= 16'hFFFF;
rommem[15170] <= 16'hFFFF;
rommem[15171] <= 16'hFFFF;
rommem[15172] <= 16'hFFFF;
rommem[15173] <= 16'hFFFF;
rommem[15174] <= 16'hFFFF;
rommem[15175] <= 16'hFFFF;
rommem[15176] <= 16'hFFFF;
rommem[15177] <= 16'hFFFF;
rommem[15178] <= 16'hFFFF;
rommem[15179] <= 16'hFFFF;
rommem[15180] <= 16'hFFFF;
rommem[15181] <= 16'hFFFF;
rommem[15182] <= 16'hFFFF;
rommem[15183] <= 16'hFFFF;
rommem[15184] <= 16'hFFFF;
rommem[15185] <= 16'hFFFF;
rommem[15186] <= 16'hFFFF;
rommem[15187] <= 16'hFFFF;
rommem[15188] <= 16'hFFFF;
rommem[15189] <= 16'hFFFF;
rommem[15190] <= 16'hFFFF;
rommem[15191] <= 16'hFFFF;
rommem[15192] <= 16'hFFFF;
rommem[15193] <= 16'hFFFF;
rommem[15194] <= 16'hFFFF;
rommem[15195] <= 16'hFFFF;
rommem[15196] <= 16'hFFFF;
rommem[15197] <= 16'hFFFF;
rommem[15198] <= 16'hFFFF;
rommem[15199] <= 16'hFFFF;
rommem[15200] <= 16'hFFFF;
rommem[15201] <= 16'hFFFF;
rommem[15202] <= 16'hFFFF;
rommem[15203] <= 16'hFFFF;
rommem[15204] <= 16'hFFFF;
rommem[15205] <= 16'hFFFF;
rommem[15206] <= 16'hFFFF;
rommem[15207] <= 16'hFFFF;
rommem[15208] <= 16'hFFFF;
rommem[15209] <= 16'hFFFF;
rommem[15210] <= 16'hFFFF;
rommem[15211] <= 16'hFFFF;
rommem[15212] <= 16'hFFFF;
rommem[15213] <= 16'hFFFF;
rommem[15214] <= 16'hFFFF;
rommem[15215] <= 16'hFFFF;
rommem[15216] <= 16'hFFFF;
rommem[15217] <= 16'hFFFF;
rommem[15218] <= 16'hFFFF;
rommem[15219] <= 16'hFFFF;
rommem[15220] <= 16'hFFFF;
rommem[15221] <= 16'hFFFF;
rommem[15222] <= 16'hFFFF;
rommem[15223] <= 16'hFFFF;
rommem[15224] <= 16'hFFFF;
rommem[15225] <= 16'hFFFF;
rommem[15226] <= 16'hFFFF;
rommem[15227] <= 16'hFFFF;
rommem[15228] <= 16'hFFFF;
rommem[15229] <= 16'hFFFF;
rommem[15230] <= 16'hFFFF;
rommem[15231] <= 16'hFFFF;
rommem[15232] <= 16'hFFFF;
rommem[15233] <= 16'hFFFF;
rommem[15234] <= 16'hFFFF;
rommem[15235] <= 16'hFFFF;
rommem[15236] <= 16'hFFFF;
rommem[15237] <= 16'hFFFF;
rommem[15238] <= 16'hFFFF;
rommem[15239] <= 16'hFFFF;
rommem[15240] <= 16'hFFFF;
rommem[15241] <= 16'hFFFF;
rommem[15242] <= 16'hFFFF;
rommem[15243] <= 16'hFFFF;
rommem[15244] <= 16'hFFFF;
rommem[15245] <= 16'hFFFF;
rommem[15246] <= 16'hFFFF;
rommem[15247] <= 16'hFFFF;
rommem[15248] <= 16'hFFFF;
rommem[15249] <= 16'hFFFF;
rommem[15250] <= 16'hFFFF;
rommem[15251] <= 16'hFFFF;
rommem[15252] <= 16'hFFFF;
rommem[15253] <= 16'hFFFF;
rommem[15254] <= 16'hFFFF;
rommem[15255] <= 16'hFFFF;
rommem[15256] <= 16'hFFFF;
rommem[15257] <= 16'hFFFF;
rommem[15258] <= 16'hFFFF;
rommem[15259] <= 16'hFFFF;
rommem[15260] <= 16'hFFFF;
rommem[15261] <= 16'hFFFF;
rommem[15262] <= 16'hFFFF;
rommem[15263] <= 16'hFFFF;
rommem[15264] <= 16'hFFFF;
rommem[15265] <= 16'hFFFF;
rommem[15266] <= 16'hFFFF;
rommem[15267] <= 16'hFFFF;
rommem[15268] <= 16'hFFFF;
rommem[15269] <= 16'hFFFF;
rommem[15270] <= 16'hFFFF;
rommem[15271] <= 16'hFFFF;
rommem[15272] <= 16'hFFFF;
rommem[15273] <= 16'hFFFF;
rommem[15274] <= 16'hFFFF;
rommem[15275] <= 16'hFFFF;
rommem[15276] <= 16'hFFFF;
rommem[15277] <= 16'hFFFF;
rommem[15278] <= 16'hFFFF;
rommem[15279] <= 16'hFFFF;
rommem[15280] <= 16'hFFFF;
rommem[15281] <= 16'hFFFF;
rommem[15282] <= 16'hFFFF;
rommem[15283] <= 16'hFFFF;
rommem[15284] <= 16'hFFFF;
rommem[15285] <= 16'hFFFF;
rommem[15286] <= 16'hFFFF;
rommem[15287] <= 16'hFFFF;
rommem[15288] <= 16'hFFFF;
rommem[15289] <= 16'hFFFF;
rommem[15290] <= 16'hFFFF;
rommem[15291] <= 16'hFFFF;
rommem[15292] <= 16'hFFFF;
rommem[15293] <= 16'hFFFF;
rommem[15294] <= 16'hFFFF;
rommem[15295] <= 16'hFFFF;
rommem[15296] <= 16'hFFFF;
rommem[15297] <= 16'hFFFF;
rommem[15298] <= 16'hFFFF;
rommem[15299] <= 16'hFFFF;
rommem[15300] <= 16'hFFFF;
rommem[15301] <= 16'hFFFF;
rommem[15302] <= 16'hFFFF;
rommem[15303] <= 16'hFFFF;
rommem[15304] <= 16'hFFFF;
rommem[15305] <= 16'hFFFF;
rommem[15306] <= 16'hFFFF;
rommem[15307] <= 16'hFFFF;
rommem[15308] <= 16'hFFFF;
rommem[15309] <= 16'hFFFF;
rommem[15310] <= 16'hFFFF;
rommem[15311] <= 16'hFFFF;
rommem[15312] <= 16'hFFFF;
rommem[15313] <= 16'hFFFF;
rommem[15314] <= 16'hFFFF;
rommem[15315] <= 16'hFFFF;
rommem[15316] <= 16'hFFFF;
rommem[15317] <= 16'hFFFF;
rommem[15318] <= 16'hFFFF;
rommem[15319] <= 16'hFFFF;
rommem[15320] <= 16'hFFFF;
rommem[15321] <= 16'hFFFF;
rommem[15322] <= 16'hFFFF;
rommem[15323] <= 16'hFFFF;
rommem[15324] <= 16'hFFFF;
rommem[15325] <= 16'hFFFF;
rommem[15326] <= 16'hFFFF;
rommem[15327] <= 16'hFFFF;
rommem[15328] <= 16'hFFFF;
rommem[15329] <= 16'hFFFF;
rommem[15330] <= 16'hFFFF;
rommem[15331] <= 16'hFFFF;
rommem[15332] <= 16'hFFFF;
rommem[15333] <= 16'hFFFF;
rommem[15334] <= 16'hFFFF;
rommem[15335] <= 16'hFFFF;
rommem[15336] <= 16'hFFFF;
rommem[15337] <= 16'hFFFF;
rommem[15338] <= 16'hFFFF;
rommem[15339] <= 16'hFFFF;
rommem[15340] <= 16'hFFFF;
rommem[15341] <= 16'hFFFF;
rommem[15342] <= 16'hFFFF;
rommem[15343] <= 16'hFFFF;
rommem[15344] <= 16'hFFFF;
rommem[15345] <= 16'hFFFF;
rommem[15346] <= 16'hFFFF;
rommem[15347] <= 16'hFFFF;
rommem[15348] <= 16'hFFFF;
rommem[15349] <= 16'hFFFF;
rommem[15350] <= 16'hFFFF;
rommem[15351] <= 16'hFFFF;
rommem[15352] <= 16'hFFFF;
rommem[15353] <= 16'hFFFF;
rommem[15354] <= 16'hFFFF;
rommem[15355] <= 16'hFFFF;
rommem[15356] <= 16'hFFFF;
rommem[15357] <= 16'hFFFF;
rommem[15358] <= 16'hFFFF;
rommem[15359] <= 16'hFFFF;
rommem[15360] <= 16'hFFFF;
rommem[15361] <= 16'hFFFF;
rommem[15362] <= 16'hFFFF;
rommem[15363] <= 16'hFFFF;
rommem[15364] <= 16'hFFFF;
rommem[15365] <= 16'hFFFF;
rommem[15366] <= 16'hFFFF;
rommem[15367] <= 16'hFFFF;
rommem[15368] <= 16'hFFFF;
rommem[15369] <= 16'hFFFF;
rommem[15370] <= 16'hFFFF;
rommem[15371] <= 16'hFFFF;
rommem[15372] <= 16'hFFFF;
rommem[15373] <= 16'hFFFF;
rommem[15374] <= 16'hFFFF;
rommem[15375] <= 16'hFFFF;
rommem[15376] <= 16'hFFFF;
rommem[15377] <= 16'hFFFF;
rommem[15378] <= 16'hFFFF;
rommem[15379] <= 16'hFFFF;
rommem[15380] <= 16'hFFFF;
rommem[15381] <= 16'hFFFF;
rommem[15382] <= 16'hFFFF;
rommem[15383] <= 16'hFFFF;
rommem[15384] <= 16'hFFFF;
rommem[15385] <= 16'hFFFF;
rommem[15386] <= 16'hFFFF;
rommem[15387] <= 16'hFFFF;
rommem[15388] <= 16'hFFFF;
rommem[15389] <= 16'hFFFF;
rommem[15390] <= 16'hFFFF;
rommem[15391] <= 16'hFFFF;
rommem[15392] <= 16'hFFFF;
rommem[15393] <= 16'hFFFF;
rommem[15394] <= 16'hFFFF;
rommem[15395] <= 16'hFFFF;
rommem[15396] <= 16'hFFFF;
rommem[15397] <= 16'hFFFF;
rommem[15398] <= 16'hFFFF;
rommem[15399] <= 16'hFFFF;
rommem[15400] <= 16'hFFFF;
rommem[15401] <= 16'hFFFF;
rommem[15402] <= 16'hFFFF;
rommem[15403] <= 16'hFFFF;
rommem[15404] <= 16'hFFFF;
rommem[15405] <= 16'hFFFF;
rommem[15406] <= 16'hFFFF;
rommem[15407] <= 16'hFFFF;
rommem[15408] <= 16'hFFFF;
rommem[15409] <= 16'hFFFF;
rommem[15410] <= 16'hFFFF;
rommem[15411] <= 16'hFFFF;
rommem[15412] <= 16'hFFFF;
rommem[15413] <= 16'hFFFF;
rommem[15414] <= 16'hFFFF;
rommem[15415] <= 16'hFFFF;
rommem[15416] <= 16'hFFFF;
rommem[15417] <= 16'hFFFF;
rommem[15418] <= 16'hFFFF;
rommem[15419] <= 16'hFFFF;
rommem[15420] <= 16'hFFFF;
rommem[15421] <= 16'hFFFF;
rommem[15422] <= 16'hFFFF;
rommem[15423] <= 16'hFFFF;
rommem[15424] <= 16'hFFFF;
rommem[15425] <= 16'hFFFF;
rommem[15426] <= 16'hFFFF;
rommem[15427] <= 16'hFFFF;
rommem[15428] <= 16'hFFFF;
rommem[15429] <= 16'hFFFF;
rommem[15430] <= 16'hFFFF;
rommem[15431] <= 16'hFFFF;
rommem[15432] <= 16'hFFFF;
rommem[15433] <= 16'hFFFF;
rommem[15434] <= 16'hFFFF;
rommem[15435] <= 16'hFFFF;
rommem[15436] <= 16'hFFFF;
rommem[15437] <= 16'hFFFF;
rommem[15438] <= 16'hFFFF;
rommem[15439] <= 16'hFFFF;
rommem[15440] <= 16'hFFFF;
rommem[15441] <= 16'hFFFF;
rommem[15442] <= 16'hFFFF;
rommem[15443] <= 16'hFFFF;
rommem[15444] <= 16'hFFFF;
rommem[15445] <= 16'hFFFF;
rommem[15446] <= 16'hFFFF;
rommem[15447] <= 16'hFFFF;
rommem[15448] <= 16'hFFFF;
rommem[15449] <= 16'hFFFF;
rommem[15450] <= 16'hFFFF;
rommem[15451] <= 16'hFFFF;
rommem[15452] <= 16'hFFFF;
rommem[15453] <= 16'hFFFF;
rommem[15454] <= 16'hFFFF;
rommem[15455] <= 16'hFFFF;
rommem[15456] <= 16'hFFFF;
rommem[15457] <= 16'hFFFF;
rommem[15458] <= 16'hFFFF;
rommem[15459] <= 16'hFFFF;
rommem[15460] <= 16'hFFFF;
rommem[15461] <= 16'hFFFF;
rommem[15462] <= 16'hFFFF;
rommem[15463] <= 16'hFFFF;
rommem[15464] <= 16'hFFFF;
rommem[15465] <= 16'hFFFF;
rommem[15466] <= 16'hFFFF;
rommem[15467] <= 16'hFFFF;
rommem[15468] <= 16'hFFFF;
rommem[15469] <= 16'hFFFF;
rommem[15470] <= 16'hFFFF;
rommem[15471] <= 16'hFFFF;
rommem[15472] <= 16'hFFFF;
rommem[15473] <= 16'hFFFF;
rommem[15474] <= 16'hFFFF;
rommem[15475] <= 16'hFFFF;
rommem[15476] <= 16'hFFFF;
rommem[15477] <= 16'hFFFF;
rommem[15478] <= 16'hFFFF;
rommem[15479] <= 16'hFFFF;
rommem[15480] <= 16'hFFFF;
rommem[15481] <= 16'hFFFF;
rommem[15482] <= 16'hFFFF;
rommem[15483] <= 16'hFFFF;
rommem[15484] <= 16'hFFFF;
rommem[15485] <= 16'hFFFF;
rommem[15486] <= 16'hFFFF;
rommem[15487] <= 16'hFFFF;
rommem[15488] <= 16'hFFFF;
rommem[15489] <= 16'hFFFF;
rommem[15490] <= 16'hFFFF;
rommem[15491] <= 16'hFFFF;
rommem[15492] <= 16'hFFFF;
rommem[15493] <= 16'hFFFF;
rommem[15494] <= 16'hFFFF;
rommem[15495] <= 16'hFFFF;
rommem[15496] <= 16'hFFFF;
rommem[15497] <= 16'hFFFF;
rommem[15498] <= 16'hFFFF;
rommem[15499] <= 16'hFFFF;
rommem[15500] <= 16'hFFFF;
rommem[15501] <= 16'hFFFF;
rommem[15502] <= 16'hFFFF;
rommem[15503] <= 16'hFFFF;
rommem[15504] <= 16'hFFFF;
rommem[15505] <= 16'hFFFF;
rommem[15506] <= 16'hFFFF;
rommem[15507] <= 16'hFFFF;
rommem[15508] <= 16'hFFFF;
rommem[15509] <= 16'hFFFF;
rommem[15510] <= 16'hFFFF;
rommem[15511] <= 16'hFFFF;
rommem[15512] <= 16'hFFFF;
rommem[15513] <= 16'hFFFF;
rommem[15514] <= 16'hFFFF;
rommem[15515] <= 16'hFFFF;
rommem[15516] <= 16'hFFFF;
rommem[15517] <= 16'hFFFF;
rommem[15518] <= 16'hFFFF;
rommem[15519] <= 16'hFFFF;
rommem[15520] <= 16'hFFFF;
rommem[15521] <= 16'hFFFF;
rommem[15522] <= 16'hFFFF;
rommem[15523] <= 16'hFFFF;
rommem[15524] <= 16'hFFFF;
rommem[15525] <= 16'hFFFF;
rommem[15526] <= 16'hFFFF;
rommem[15527] <= 16'hFFFF;
rommem[15528] <= 16'hFFFF;
rommem[15529] <= 16'hFFFF;
rommem[15530] <= 16'hFFFF;
rommem[15531] <= 16'hFFFF;
rommem[15532] <= 16'hFFFF;
rommem[15533] <= 16'hFFFF;
rommem[15534] <= 16'hFFFF;
rommem[15535] <= 16'hFFFF;
rommem[15536] <= 16'hFFFF;
rommem[15537] <= 16'hFFFF;
rommem[15538] <= 16'hFFFF;
rommem[15539] <= 16'hFFFF;
rommem[15540] <= 16'hFFFF;
rommem[15541] <= 16'hFFFF;
rommem[15542] <= 16'hFFFF;
rommem[15543] <= 16'hFFFF;
rommem[15544] <= 16'hFFFF;
rommem[15545] <= 16'hFFFF;
rommem[15546] <= 16'hFFFF;
rommem[15547] <= 16'hFFFF;
rommem[15548] <= 16'hFFFF;
rommem[15549] <= 16'hFFFF;
rommem[15550] <= 16'hFFFF;
rommem[15551] <= 16'hFFFF;
rommem[15552] <= 16'hFFFF;
rommem[15553] <= 16'hFFFF;
rommem[15554] <= 16'hFFFF;
rommem[15555] <= 16'hFFFF;
rommem[15556] <= 16'hFFFF;
rommem[15557] <= 16'hFFFF;
rommem[15558] <= 16'hFFFF;
rommem[15559] <= 16'hFFFF;
rommem[15560] <= 16'hFFFF;
rommem[15561] <= 16'hFFFF;
rommem[15562] <= 16'hFFFF;
rommem[15563] <= 16'hFFFF;
rommem[15564] <= 16'hFFFF;
rommem[15565] <= 16'hFFFF;
rommem[15566] <= 16'hFFFF;
rommem[15567] <= 16'hFFFF;
rommem[15568] <= 16'hFFFF;
rommem[15569] <= 16'hFFFF;
rommem[15570] <= 16'hFFFF;
rommem[15571] <= 16'hFFFF;
rommem[15572] <= 16'hFFFF;
rommem[15573] <= 16'hFFFF;
rommem[15574] <= 16'hFFFF;
rommem[15575] <= 16'hFFFF;
rommem[15576] <= 16'hFFFF;
rommem[15577] <= 16'hFFFF;
rommem[15578] <= 16'hFFFF;
rommem[15579] <= 16'hFFFF;
rommem[15580] <= 16'hFFFF;
rommem[15581] <= 16'hFFFF;
rommem[15582] <= 16'hFFFF;
rommem[15583] <= 16'hFFFF;
rommem[15584] <= 16'hFFFF;
rommem[15585] <= 16'hFFFF;
rommem[15586] <= 16'hFFFF;
rommem[15587] <= 16'hFFFF;
rommem[15588] <= 16'hFFFF;
rommem[15589] <= 16'hFFFF;
rommem[15590] <= 16'hFFFF;
rommem[15591] <= 16'hFFFF;
rommem[15592] <= 16'hFFFF;
rommem[15593] <= 16'hFFFF;
rommem[15594] <= 16'hFFFF;
rommem[15595] <= 16'hFFFF;
rommem[15596] <= 16'hFFFF;
rommem[15597] <= 16'hFFFF;
rommem[15598] <= 16'hFFFF;
rommem[15599] <= 16'hFFFF;
rommem[15600] <= 16'hFFFF;
rommem[15601] <= 16'hFFFF;
rommem[15602] <= 16'hFFFF;
rommem[15603] <= 16'hFFFF;
rommem[15604] <= 16'hFFFF;
rommem[15605] <= 16'hFFFF;
rommem[15606] <= 16'hFFFF;
rommem[15607] <= 16'hFFFF;
rommem[15608] <= 16'hFFFF;
rommem[15609] <= 16'hFFFF;
rommem[15610] <= 16'hFFFF;
rommem[15611] <= 16'hFFFF;
rommem[15612] <= 16'hFFFF;
rommem[15613] <= 16'hFFFF;
rommem[15614] <= 16'hFFFF;
rommem[15615] <= 16'hFFFF;
rommem[15616] <= 16'hFFFF;
rommem[15617] <= 16'hFFFF;
rommem[15618] <= 16'hFFFF;
rommem[15619] <= 16'hFFFF;
rommem[15620] <= 16'hFFFF;
rommem[15621] <= 16'hFFFF;
rommem[15622] <= 16'hFFFF;
rommem[15623] <= 16'hFFFF;
rommem[15624] <= 16'hFFFF;
rommem[15625] <= 16'hFFFF;
rommem[15626] <= 16'hFFFF;
rommem[15627] <= 16'hFFFF;
rommem[15628] <= 16'hFFFF;
rommem[15629] <= 16'hFFFF;
rommem[15630] <= 16'hFFFF;
rommem[15631] <= 16'hFFFF;
rommem[15632] <= 16'hFFFF;
rommem[15633] <= 16'hFFFF;
rommem[15634] <= 16'hFFFF;
rommem[15635] <= 16'hFFFF;
rommem[15636] <= 16'hFFFF;
rommem[15637] <= 16'hFFFF;
rommem[15638] <= 16'hFFFF;
rommem[15639] <= 16'hFFFF;
rommem[15640] <= 16'hFFFF;
rommem[15641] <= 16'hFFFF;
rommem[15642] <= 16'hFFFF;
rommem[15643] <= 16'hFFFF;
rommem[15644] <= 16'hFFFF;
rommem[15645] <= 16'hFFFF;
rommem[15646] <= 16'hFFFF;
rommem[15647] <= 16'hFFFF;
rommem[15648] <= 16'hFFFF;
rommem[15649] <= 16'hFFFF;
rommem[15650] <= 16'hFFFF;
rommem[15651] <= 16'hFFFF;
rommem[15652] <= 16'hFFFF;
rommem[15653] <= 16'hFFFF;
rommem[15654] <= 16'hFFFF;
rommem[15655] <= 16'hFFFF;
rommem[15656] <= 16'hFFFF;
rommem[15657] <= 16'hFFFF;
rommem[15658] <= 16'hFFFF;
rommem[15659] <= 16'hFFFF;
rommem[15660] <= 16'hFFFF;
rommem[15661] <= 16'hFFFF;
rommem[15662] <= 16'hFFFF;
rommem[15663] <= 16'hFFFF;
rommem[15664] <= 16'hFFFF;
rommem[15665] <= 16'hFFFF;
rommem[15666] <= 16'hFFFF;
rommem[15667] <= 16'hFFFF;
rommem[15668] <= 16'hFFFF;
rommem[15669] <= 16'hFFFF;
rommem[15670] <= 16'hFFFF;
rommem[15671] <= 16'hFFFF;
rommem[15672] <= 16'hFFFF;
rommem[15673] <= 16'hFFFF;
rommem[15674] <= 16'hFFFF;
rommem[15675] <= 16'hFFFF;
rommem[15676] <= 16'hFFFF;
rommem[15677] <= 16'hFFFF;
rommem[15678] <= 16'hFFFF;
rommem[15679] <= 16'hFFFF;
rommem[15680] <= 16'hFFFF;
rommem[15681] <= 16'hFFFF;
rommem[15682] <= 16'hFFFF;
rommem[15683] <= 16'hFFFF;
rommem[15684] <= 16'hFFFF;
rommem[15685] <= 16'hFFFF;
rommem[15686] <= 16'hFFFF;
rommem[15687] <= 16'hFFFF;
rommem[15688] <= 16'hFFFF;
rommem[15689] <= 16'hFFFF;
rommem[15690] <= 16'hFFFF;
rommem[15691] <= 16'hFFFF;
rommem[15692] <= 16'hFFFF;
rommem[15693] <= 16'hFFFF;
rommem[15694] <= 16'hFFFF;
rommem[15695] <= 16'hFFFF;
rommem[15696] <= 16'hFFFF;
rommem[15697] <= 16'hFFFF;
rommem[15698] <= 16'hFFFF;
rommem[15699] <= 16'hFFFF;
rommem[15700] <= 16'hFFFF;
rommem[15701] <= 16'hFFFF;
rommem[15702] <= 16'hFFFF;
rommem[15703] <= 16'hFFFF;
rommem[15704] <= 16'hFFFF;
rommem[15705] <= 16'hFFFF;
rommem[15706] <= 16'hFFFF;
rommem[15707] <= 16'hFFFF;
rommem[15708] <= 16'hFFFF;
rommem[15709] <= 16'hFFFF;
rommem[15710] <= 16'hFFFF;
rommem[15711] <= 16'hFFFF;
rommem[15712] <= 16'hFFFF;
rommem[15713] <= 16'hFFFF;
rommem[15714] <= 16'hFFFF;
rommem[15715] <= 16'hFFFF;
rommem[15716] <= 16'hFFFF;
rommem[15717] <= 16'hFFFF;
rommem[15718] <= 16'hFFFF;
rommem[15719] <= 16'hFFFF;
rommem[15720] <= 16'hFFFF;
rommem[15721] <= 16'hFFFF;
rommem[15722] <= 16'hFFFF;
rommem[15723] <= 16'hFFFF;
rommem[15724] <= 16'hFFFF;
rommem[15725] <= 16'hFFFF;
rommem[15726] <= 16'hFFFF;
rommem[15727] <= 16'hFFFF;
rommem[15728] <= 16'hFFFF;
rommem[15729] <= 16'hFFFF;
rommem[15730] <= 16'hFFFF;
rommem[15731] <= 16'hFFFF;
rommem[15732] <= 16'hFFFF;
rommem[15733] <= 16'hFFFF;
rommem[15734] <= 16'hFFFF;
rommem[15735] <= 16'hFFFF;
rommem[15736] <= 16'hFFFF;
rommem[15737] <= 16'hFFFF;
rommem[15738] <= 16'hFFFF;
rommem[15739] <= 16'hFFFF;
rommem[15740] <= 16'hFFFF;
rommem[15741] <= 16'hFFFF;
rommem[15742] <= 16'hFFFF;
rommem[15743] <= 16'hFFFF;
rommem[15744] <= 16'hFFFF;
rommem[15745] <= 16'hFFFF;
rommem[15746] <= 16'hFFFF;
rommem[15747] <= 16'hFFFF;
rommem[15748] <= 16'hFFFF;
rommem[15749] <= 16'hFFFF;
rommem[15750] <= 16'hFFFF;
rommem[15751] <= 16'hFFFF;
rommem[15752] <= 16'hFFFF;
rommem[15753] <= 16'hFFFF;
rommem[15754] <= 16'hFFFF;
rommem[15755] <= 16'hFFFF;
rommem[15756] <= 16'hFFFF;
rommem[15757] <= 16'hFFFF;
rommem[15758] <= 16'hFFFF;
rommem[15759] <= 16'hFFFF;
rommem[15760] <= 16'hFFFF;
rommem[15761] <= 16'hFFFF;
rommem[15762] <= 16'hFFFF;
rommem[15763] <= 16'hFFFF;
rommem[15764] <= 16'hFFFF;
rommem[15765] <= 16'hFFFF;
rommem[15766] <= 16'hFFFF;
rommem[15767] <= 16'hFFFF;
rommem[15768] <= 16'hFFFF;
rommem[15769] <= 16'hFFFF;
rommem[15770] <= 16'hFFFF;
rommem[15771] <= 16'hFFFF;
rommem[15772] <= 16'hFFFF;
rommem[15773] <= 16'hFFFF;
rommem[15774] <= 16'hFFFF;
rommem[15775] <= 16'hFFFF;
rommem[15776] <= 16'hFFFF;
rommem[15777] <= 16'hFFFF;
rommem[15778] <= 16'hFFFF;
rommem[15779] <= 16'hFFFF;
rommem[15780] <= 16'hFFFF;
rommem[15781] <= 16'hFFFF;
rommem[15782] <= 16'hFFFF;
rommem[15783] <= 16'hFFFF;
rommem[15784] <= 16'hFFFF;
rommem[15785] <= 16'hFFFF;
rommem[15786] <= 16'hFFFF;
rommem[15787] <= 16'hFFFF;
rommem[15788] <= 16'hFFFF;
rommem[15789] <= 16'hFFFF;
rommem[15790] <= 16'hFFFF;
rommem[15791] <= 16'hFFFF;
rommem[15792] <= 16'hFFFF;
rommem[15793] <= 16'hFFFF;
rommem[15794] <= 16'hFFFF;
rommem[15795] <= 16'hFFFF;
rommem[15796] <= 16'hFFFF;
rommem[15797] <= 16'hFFFF;
rommem[15798] <= 16'hFFFF;
rommem[15799] <= 16'hFFFF;
rommem[15800] <= 16'hFFFF;
rommem[15801] <= 16'hFFFF;
rommem[15802] <= 16'hFFFF;
rommem[15803] <= 16'hFFFF;
rommem[15804] <= 16'hFFFF;
rommem[15805] <= 16'hFFFF;
rommem[15806] <= 16'hFFFF;
rommem[15807] <= 16'hFFFF;
rommem[15808] <= 16'hFFFF;
rommem[15809] <= 16'hFFFF;
rommem[15810] <= 16'hFFFF;
rommem[15811] <= 16'hFFFF;
rommem[15812] <= 16'hFFFF;
rommem[15813] <= 16'hFFFF;
rommem[15814] <= 16'hFFFF;
rommem[15815] <= 16'hFFFF;
rommem[15816] <= 16'hFFFF;
rommem[15817] <= 16'hFFFF;
rommem[15818] <= 16'hFFFF;
rommem[15819] <= 16'hFFFF;
rommem[15820] <= 16'hFFFF;
rommem[15821] <= 16'hFFFF;
rommem[15822] <= 16'hFFFF;
rommem[15823] <= 16'hFFFF;
rommem[15824] <= 16'hFFFF;
rommem[15825] <= 16'hFFFF;
rommem[15826] <= 16'hFFFF;
rommem[15827] <= 16'hFFFF;
rommem[15828] <= 16'hFFFF;
rommem[15829] <= 16'hFFFF;
rommem[15830] <= 16'hFFFF;
rommem[15831] <= 16'hFFFF;
rommem[15832] <= 16'hFFFF;
rommem[15833] <= 16'hFFFF;
rommem[15834] <= 16'hFFFF;
rommem[15835] <= 16'hFFFF;
rommem[15836] <= 16'hFFFF;
rommem[15837] <= 16'hFFFF;
rommem[15838] <= 16'hFFFF;
rommem[15839] <= 16'hFFFF;
rommem[15840] <= 16'hFFFF;
rommem[15841] <= 16'hFFFF;
rommem[15842] <= 16'hFFFF;
rommem[15843] <= 16'hFFFF;
rommem[15844] <= 16'hFFFF;
rommem[15845] <= 16'hFFFF;
rommem[15846] <= 16'hFFFF;
rommem[15847] <= 16'hFFFF;
rommem[15848] <= 16'hFFFF;
rommem[15849] <= 16'hFFFF;
rommem[15850] <= 16'hFFFF;
rommem[15851] <= 16'hFFFF;
rommem[15852] <= 16'hFFFF;
rommem[15853] <= 16'hFFFF;
rommem[15854] <= 16'hFFFF;
rommem[15855] <= 16'hFFFF;
rommem[15856] <= 16'hFFFF;
rommem[15857] <= 16'hFFFF;
rommem[15858] <= 16'hFFFF;
rommem[15859] <= 16'hFFFF;
rommem[15860] <= 16'hFFFF;
rommem[15861] <= 16'hFFFF;
rommem[15862] <= 16'hFFFF;
rommem[15863] <= 16'hFFFF;
rommem[15864] <= 16'hFFFF;
rommem[15865] <= 16'hFFFF;
rommem[15866] <= 16'hFFFF;
rommem[15867] <= 16'hFFFF;
rommem[15868] <= 16'hFFFF;
rommem[15869] <= 16'hFFFF;
rommem[15870] <= 16'hFFFF;
rommem[15871] <= 16'hFFFF;
rommem[15872] <= 16'hFFFF;
rommem[15873] <= 16'hFFFF;
rommem[15874] <= 16'hFFFF;
rommem[15875] <= 16'hFFFF;
rommem[15876] <= 16'hFFFF;
rommem[15877] <= 16'hFFFF;
rommem[15878] <= 16'hFFFF;
rommem[15879] <= 16'hFFFF;
rommem[15880] <= 16'hFFFF;
rommem[15881] <= 16'hFFFF;
rommem[15882] <= 16'hFFFF;
rommem[15883] <= 16'hFFFF;
rommem[15884] <= 16'hFFFF;
rommem[15885] <= 16'hFFFF;
rommem[15886] <= 16'hFFFF;
rommem[15887] <= 16'hFFFF;
rommem[15888] <= 16'hFFFF;
rommem[15889] <= 16'hFFFF;
rommem[15890] <= 16'hFFFF;
rommem[15891] <= 16'hFFFF;
rommem[15892] <= 16'hFFFF;
rommem[15893] <= 16'hFFFF;
rommem[15894] <= 16'hFFFF;
rommem[15895] <= 16'hFFFF;
rommem[15896] <= 16'hFFFF;
rommem[15897] <= 16'hFFFF;
rommem[15898] <= 16'hFFFF;
rommem[15899] <= 16'hFFFF;
rommem[15900] <= 16'hFFFF;
rommem[15901] <= 16'hFFFF;
rommem[15902] <= 16'hFFFF;
rommem[15903] <= 16'hFFFF;
rommem[15904] <= 16'hFFFF;
rommem[15905] <= 16'hFFFF;
rommem[15906] <= 16'hFFFF;
rommem[15907] <= 16'hFFFF;
rommem[15908] <= 16'hFFFF;
rommem[15909] <= 16'hFFFF;
rommem[15910] <= 16'hFFFF;
rommem[15911] <= 16'hFFFF;
rommem[15912] <= 16'hFFFF;
rommem[15913] <= 16'hFFFF;
rommem[15914] <= 16'hFFFF;
rommem[15915] <= 16'hFFFF;
rommem[15916] <= 16'hFFFF;
rommem[15917] <= 16'hFFFF;
rommem[15918] <= 16'hFFFF;
rommem[15919] <= 16'hFFFF;
rommem[15920] <= 16'hFFFF;
rommem[15921] <= 16'hFFFF;
rommem[15922] <= 16'hFFFF;
rommem[15923] <= 16'hFFFF;
rommem[15924] <= 16'hFFFF;
rommem[15925] <= 16'hFFFF;
rommem[15926] <= 16'hFFFF;
rommem[15927] <= 16'hFFFF;
rommem[15928] <= 16'hFFFF;
rommem[15929] <= 16'hFFFF;
rommem[15930] <= 16'hFFFF;
rommem[15931] <= 16'hFFFF;
rommem[15932] <= 16'hFFFF;
rommem[15933] <= 16'hFFFF;
rommem[15934] <= 16'hFFFF;
rommem[15935] <= 16'hFFFF;
rommem[15936] <= 16'hFFFF;
rommem[15937] <= 16'hFFFF;
rommem[15938] <= 16'hFFFF;
rommem[15939] <= 16'hFFFF;
rommem[15940] <= 16'hFFFF;
rommem[15941] <= 16'hFFFF;
rommem[15942] <= 16'hFFFF;
rommem[15943] <= 16'hFFFF;
rommem[15944] <= 16'hFFFF;
rommem[15945] <= 16'hFFFF;
rommem[15946] <= 16'hFFFF;
rommem[15947] <= 16'hFFFF;
rommem[15948] <= 16'hFFFF;
rommem[15949] <= 16'hFFFF;
rommem[15950] <= 16'hFFFF;
rommem[15951] <= 16'hFFFF;
rommem[15952] <= 16'hFFFF;
rommem[15953] <= 16'hFFFF;
rommem[15954] <= 16'hFFFF;
rommem[15955] <= 16'hFFFF;
rommem[15956] <= 16'hFFFF;
rommem[15957] <= 16'hFFFF;
rommem[15958] <= 16'hFFFF;
rommem[15959] <= 16'hFFFF;
rommem[15960] <= 16'hFFFF;
rommem[15961] <= 16'hFFFF;
rommem[15962] <= 16'hFFFF;
rommem[15963] <= 16'hFFFF;
rommem[15964] <= 16'hFFFF;
rommem[15965] <= 16'hFFFF;
rommem[15966] <= 16'hFFFF;
rommem[15967] <= 16'hFFFF;
rommem[15968] <= 16'hFFFF;
rommem[15969] <= 16'hFFFF;
rommem[15970] <= 16'hFFFF;
rommem[15971] <= 16'hFFFF;
rommem[15972] <= 16'hFFFF;
rommem[15973] <= 16'hFFFF;
rommem[15974] <= 16'hFFFF;
rommem[15975] <= 16'hFFFF;
rommem[15976] <= 16'hFFFF;
rommem[15977] <= 16'hFFFF;
rommem[15978] <= 16'hFFFF;
rommem[15979] <= 16'hFFFF;
rommem[15980] <= 16'hFFFF;
rommem[15981] <= 16'hFFFF;
rommem[15982] <= 16'hFFFF;
rommem[15983] <= 16'hFFFF;
rommem[15984] <= 16'hFFFF;
rommem[15985] <= 16'hFFFF;
rommem[15986] <= 16'hFFFF;
rommem[15987] <= 16'hFFFF;
rommem[15988] <= 16'hFFFF;
rommem[15989] <= 16'hFFFF;
rommem[15990] <= 16'hFFFF;
rommem[15991] <= 16'hFFFF;
rommem[15992] <= 16'hFFFF;
rommem[15993] <= 16'hFFFF;
rommem[15994] <= 16'hFFFF;
rommem[15995] <= 16'hFFFF;
rommem[15996] <= 16'hFFFF;
rommem[15997] <= 16'hFFFF;
rommem[15998] <= 16'hFFFF;
rommem[15999] <= 16'hFFFF;
rommem[16000] <= 16'hFFFF;
rommem[16001] <= 16'hFFFF;
rommem[16002] <= 16'hFFFF;
rommem[16003] <= 16'hFFFF;
rommem[16004] <= 16'hFFFF;
rommem[16005] <= 16'hFFFF;
rommem[16006] <= 16'hFFFF;
rommem[16007] <= 16'hFFFF;
rommem[16008] <= 16'hFFFF;
rommem[16009] <= 16'hFFFF;
rommem[16010] <= 16'hFFFF;
rommem[16011] <= 16'hFFFF;
rommem[16012] <= 16'hFFFF;
rommem[16013] <= 16'hFFFF;
rommem[16014] <= 16'hFFFF;
rommem[16015] <= 16'hFFFF;
rommem[16016] <= 16'hFFFF;
rommem[16017] <= 16'hFFFF;
rommem[16018] <= 16'hFFFF;
rommem[16019] <= 16'hFFFF;
rommem[16020] <= 16'hFFFF;
rommem[16021] <= 16'hFFFF;
rommem[16022] <= 16'hFFFF;
rommem[16023] <= 16'hFFFF;
rommem[16024] <= 16'hFFFF;
rommem[16025] <= 16'hFFFF;
rommem[16026] <= 16'hFFFF;
rommem[16027] <= 16'hFFFF;
rommem[16028] <= 16'hFFFF;
rommem[16029] <= 16'hFFFF;
rommem[16030] <= 16'hFFFF;
rommem[16031] <= 16'hFFFF;
rommem[16032] <= 16'hFFFF;
rommem[16033] <= 16'hFFFF;
rommem[16034] <= 16'hFFFF;
rommem[16035] <= 16'hFFFF;
rommem[16036] <= 16'hFFFF;
rommem[16037] <= 16'hFFFF;
rommem[16038] <= 16'hFFFF;
rommem[16039] <= 16'hFFFF;
rommem[16040] <= 16'hFFFF;
rommem[16041] <= 16'hFFFF;
rommem[16042] <= 16'hFFFF;
rommem[16043] <= 16'hFFFF;
rommem[16044] <= 16'hFFFF;
rommem[16045] <= 16'hFFFF;
rommem[16046] <= 16'hFFFF;
rommem[16047] <= 16'hFFFF;
rommem[16048] <= 16'hFFFF;
rommem[16049] <= 16'hFFFF;
rommem[16050] <= 16'hFFFF;
rommem[16051] <= 16'hFFFF;
rommem[16052] <= 16'hFFFF;
rommem[16053] <= 16'hFFFF;
rommem[16054] <= 16'hFFFF;
rommem[16055] <= 16'hFFFF;
rommem[16056] <= 16'hFFFF;
rommem[16057] <= 16'hFFFF;
rommem[16058] <= 16'hFFFF;
rommem[16059] <= 16'hFFFF;
rommem[16060] <= 16'hFFFF;
rommem[16061] <= 16'hFFFF;
rommem[16062] <= 16'hFFFF;
rommem[16063] <= 16'hFFFF;
rommem[16064] <= 16'hFFFF;
rommem[16065] <= 16'hFFFF;
rommem[16066] <= 16'hFFFF;
rommem[16067] <= 16'hFFFF;
rommem[16068] <= 16'hFFFF;
rommem[16069] <= 16'hFFFF;
rommem[16070] <= 16'hFFFF;
rommem[16071] <= 16'hFFFF;
rommem[16072] <= 16'hFFFF;
rommem[16073] <= 16'hFFFF;
rommem[16074] <= 16'hFFFF;
rommem[16075] <= 16'hFFFF;
rommem[16076] <= 16'hFFFF;
rommem[16077] <= 16'hFFFF;
rommem[16078] <= 16'hFFFF;
rommem[16079] <= 16'hFFFF;
rommem[16080] <= 16'hFFFF;
rommem[16081] <= 16'hFFFF;
rommem[16082] <= 16'hFFFF;
rommem[16083] <= 16'hFFFF;
rommem[16084] <= 16'hFFFF;
rommem[16085] <= 16'hFFFF;
rommem[16086] <= 16'hFFFF;
rommem[16087] <= 16'hFFFF;
rommem[16088] <= 16'hFFFF;
rommem[16089] <= 16'hFFFF;
rommem[16090] <= 16'hFFFF;
rommem[16091] <= 16'hFFFF;
rommem[16092] <= 16'hFFFF;
rommem[16093] <= 16'hFFFF;
rommem[16094] <= 16'hFFFF;
rommem[16095] <= 16'hFFFF;
rommem[16096] <= 16'hFFFF;
rommem[16097] <= 16'hFFFF;
rommem[16098] <= 16'hFFFF;
rommem[16099] <= 16'hFFFF;
rommem[16100] <= 16'hFFFF;
rommem[16101] <= 16'hFFFF;
rommem[16102] <= 16'hFFFF;
rommem[16103] <= 16'hFFFF;
rommem[16104] <= 16'hFFFF;
rommem[16105] <= 16'hFFFF;
rommem[16106] <= 16'hFFFF;
rommem[16107] <= 16'hFFFF;
rommem[16108] <= 16'hFFFF;
rommem[16109] <= 16'hFFFF;
rommem[16110] <= 16'hFFFF;
rommem[16111] <= 16'hFFFF;
rommem[16112] <= 16'hFFFF;
rommem[16113] <= 16'hFFFF;
rommem[16114] <= 16'hFFFF;
rommem[16115] <= 16'hFFFF;
rommem[16116] <= 16'hFFFF;
rommem[16117] <= 16'hFFFF;
rommem[16118] <= 16'hFFFF;
rommem[16119] <= 16'hFFFF;
rommem[16120] <= 16'hFFFF;
rommem[16121] <= 16'hFFFF;
rommem[16122] <= 16'hFFFF;
rommem[16123] <= 16'hFFFF;
rommem[16124] <= 16'hFFFF;
rommem[16125] <= 16'hFFFF;
rommem[16126] <= 16'hFFFF;
rommem[16127] <= 16'hFFFF;
rommem[16128] <= 16'hFFFF;
rommem[16129] <= 16'hFFFF;
rommem[16130] <= 16'hFFFF;
rommem[16131] <= 16'hFFFF;
rommem[16132] <= 16'hFFFF;
rommem[16133] <= 16'hFFFF;
rommem[16134] <= 16'hFFFF;
rommem[16135] <= 16'hFFFF;
rommem[16136] <= 16'hFFFF;
rommem[16137] <= 16'hFFFF;
rommem[16138] <= 16'hFFFF;
rommem[16139] <= 16'hFFFF;
rommem[16140] <= 16'hFFFF;
rommem[16141] <= 16'hFFFF;
rommem[16142] <= 16'hFFFF;
rommem[16143] <= 16'hFFFF;
rommem[16144] <= 16'hFFFF;
rommem[16145] <= 16'hFFFF;
rommem[16146] <= 16'hFFFF;
rommem[16147] <= 16'hFFFF;
rommem[16148] <= 16'hFFFF;
rommem[16149] <= 16'hFFFF;
rommem[16150] <= 16'hFFFF;
rommem[16151] <= 16'hFFFF;
rommem[16152] <= 16'hFFFF;
rommem[16153] <= 16'hFFFF;
rommem[16154] <= 16'hFFFF;
rommem[16155] <= 16'hFFFF;
rommem[16156] <= 16'hFFFF;
rommem[16157] <= 16'hFFFF;
rommem[16158] <= 16'hFFFF;
rommem[16159] <= 16'hFFFF;
rommem[16160] <= 16'hFFFF;
rommem[16161] <= 16'hFFFF;
rommem[16162] <= 16'hFFFF;
rommem[16163] <= 16'hFFFF;
rommem[16164] <= 16'hFFFF;
rommem[16165] <= 16'hFFFF;
rommem[16166] <= 16'hFFFF;
rommem[16167] <= 16'hFFFF;
rommem[16168] <= 16'hFFFF;
rommem[16169] <= 16'hFFFF;
rommem[16170] <= 16'hFFFF;
rommem[16171] <= 16'hFFFF;
rommem[16172] <= 16'hFFFF;
rommem[16173] <= 16'hFFFF;
rommem[16174] <= 16'hFFFF;
rommem[16175] <= 16'hFFFF;
rommem[16176] <= 16'hFFFF;
rommem[16177] <= 16'hFFFF;
rommem[16178] <= 16'hFFFF;
rommem[16179] <= 16'hFFFF;
rommem[16180] <= 16'hFFFF;
rommem[16181] <= 16'hFFFF;
rommem[16182] <= 16'hFFFF;
rommem[16183] <= 16'hFFFF;
rommem[16184] <= 16'hFFFF;
rommem[16185] <= 16'hFFFF;
rommem[16186] <= 16'hFFFF;
rommem[16187] <= 16'hFFFF;
rommem[16188] <= 16'hFFFF;
rommem[16189] <= 16'hFFFF;
rommem[16190] <= 16'hFFFF;
rommem[16191] <= 16'hFFFF;
rommem[16192] <= 16'hFFFF;
rommem[16193] <= 16'hFFFF;
rommem[16194] <= 16'hFFFF;
rommem[16195] <= 16'hFFFF;
rommem[16196] <= 16'hFFFF;
rommem[16197] <= 16'hFFFF;
rommem[16198] <= 16'hFFFF;
rommem[16199] <= 16'hFFFF;
rommem[16200] <= 16'hFFFF;
rommem[16201] <= 16'hFFFF;
rommem[16202] <= 16'hFFFF;
rommem[16203] <= 16'hFFFF;
rommem[16204] <= 16'hFFFF;
rommem[16205] <= 16'hFFFF;
rommem[16206] <= 16'hFFFF;
rommem[16207] <= 16'hFFFF;
rommem[16208] <= 16'hFFFF;
rommem[16209] <= 16'hFFFF;
rommem[16210] <= 16'hFFFF;
rommem[16211] <= 16'hFFFF;
rommem[16212] <= 16'hFFFF;
rommem[16213] <= 16'hFFFF;
rommem[16214] <= 16'hFFFF;
rommem[16215] <= 16'hFFFF;
rommem[16216] <= 16'hFFFF;
rommem[16217] <= 16'hFFFF;
rommem[16218] <= 16'hFFFF;
rommem[16219] <= 16'hFFFF;
rommem[16220] <= 16'hFFFF;
rommem[16221] <= 16'hFFFF;
rommem[16222] <= 16'hFFFF;
rommem[16223] <= 16'hFFFF;
rommem[16224] <= 16'hFFFF;
rommem[16225] <= 16'hFFFF;
rommem[16226] <= 16'hFFFF;
rommem[16227] <= 16'hFFFF;
rommem[16228] <= 16'hFFFF;
rommem[16229] <= 16'hFFFF;
rommem[16230] <= 16'hFFFF;
rommem[16231] <= 16'hFFFF;
rommem[16232] <= 16'hFFFF;
rommem[16233] <= 16'hFFFF;
rommem[16234] <= 16'hFFFF;
rommem[16235] <= 16'hFFFF;
rommem[16236] <= 16'hFFFF;
rommem[16237] <= 16'hFFFF;
rommem[16238] <= 16'hFFFF;
rommem[16239] <= 16'hFFFF;
rommem[16240] <= 16'hFFFF;
rommem[16241] <= 16'hFFFF;
rommem[16242] <= 16'hFFFF;
rommem[16243] <= 16'hFFFF;
rommem[16244] <= 16'hFFFF;
rommem[16245] <= 16'hFFFF;
rommem[16246] <= 16'hFFFF;
rommem[16247] <= 16'hFFFF;
rommem[16248] <= 16'hFFFF;
rommem[16249] <= 16'hFFFF;
rommem[16250] <= 16'hFFFF;
rommem[16251] <= 16'hFFFF;
rommem[16252] <= 16'hFFFF;
rommem[16253] <= 16'hFFFF;
rommem[16254] <= 16'hFFFF;
rommem[16255] <= 16'hFFFF;
rommem[16256] <= 16'hFFFF;
rommem[16257] <= 16'hFFFF;
rommem[16258] <= 16'hFFFF;
rommem[16259] <= 16'hFFFF;
rommem[16260] <= 16'hFFFF;
rommem[16261] <= 16'hFFFF;
rommem[16262] <= 16'hFFFF;
rommem[16263] <= 16'hFFFF;
rommem[16264] <= 16'hFFFF;
rommem[16265] <= 16'hFFFF;
rommem[16266] <= 16'hFFFF;
rommem[16267] <= 16'hFFFF;
rommem[16268] <= 16'hFFFF;
rommem[16269] <= 16'hFFFF;
rommem[16270] <= 16'hFFFF;
rommem[16271] <= 16'hFFFF;
rommem[16272] <= 16'hFFFF;
rommem[16273] <= 16'hFFFF;
rommem[16274] <= 16'hFFFF;
rommem[16275] <= 16'hFFFF;
rommem[16276] <= 16'hFFFF;
rommem[16277] <= 16'hFFFF;
rommem[16278] <= 16'hFFFF;
rommem[16279] <= 16'hFFFF;
rommem[16280] <= 16'hFFFF;
rommem[16281] <= 16'hFFFF;
rommem[16282] <= 16'hFFFF;
rommem[16283] <= 16'hFFFF;
rommem[16284] <= 16'hFFFF;
rommem[16285] <= 16'hFFFF;
rommem[16286] <= 16'hFFFF;
rommem[16287] <= 16'hFFFF;
rommem[16288] <= 16'hFFFF;
rommem[16289] <= 16'hFFFF;
rommem[16290] <= 16'hFFFF;
rommem[16291] <= 16'hFFFF;
rommem[16292] <= 16'hFFFF;
rommem[16293] <= 16'hFFFF;
rommem[16294] <= 16'hFFFF;
rommem[16295] <= 16'hFFFF;
rommem[16296] <= 16'hFFFF;
rommem[16297] <= 16'hFFFF;
rommem[16298] <= 16'hFFFF;
rommem[16299] <= 16'hFFFF;
rommem[16300] <= 16'hFFFF;
rommem[16301] <= 16'hFFFF;
rommem[16302] <= 16'hFFFF;
rommem[16303] <= 16'hFFFF;
rommem[16304] <= 16'hFFFF;
rommem[16305] <= 16'hFFFF;
rommem[16306] <= 16'hFFFF;
rommem[16307] <= 16'hFFFF;
rommem[16308] <= 16'hFFFF;
rommem[16309] <= 16'hFFFF;
rommem[16310] <= 16'hFFFF;
rommem[16311] <= 16'hFFFF;
rommem[16312] <= 16'hFFFF;
rommem[16313] <= 16'hFFFF;
rommem[16314] <= 16'hFFFF;
rommem[16315] <= 16'hFFFF;
rommem[16316] <= 16'hFFFF;
rommem[16317] <= 16'hFFFF;
rommem[16318] <= 16'hFFFF;
rommem[16319] <= 16'hFFFF;
rommem[16320] <= 16'hFFFF;
rommem[16321] <= 16'hFFFF;
rommem[16322] <= 16'hFFFF;
rommem[16323] <= 16'hFFFF;
rommem[16324] <= 16'hFFFF;
rommem[16325] <= 16'hFFFF;
rommem[16326] <= 16'hFFFF;
rommem[16327] <= 16'hFFFF;
rommem[16328] <= 16'hFFFF;
rommem[16329] <= 16'hFFFF;
rommem[16330] <= 16'hFFFF;
rommem[16331] <= 16'hFFFF;
rommem[16332] <= 16'hFFFF;
rommem[16333] <= 16'hFFFF;
rommem[16334] <= 16'hFFFF;
rommem[16335] <= 16'hFFFF;
rommem[16336] <= 16'hFFFF;
rommem[16337] <= 16'hFFFF;
rommem[16338] <= 16'hFFFF;
rommem[16339] <= 16'hFFFF;
rommem[16340] <= 16'hFFFF;
rommem[16341] <= 16'hFFFF;
rommem[16342] <= 16'hFFFF;
rommem[16343] <= 16'hFFFF;
rommem[16344] <= 16'hFFFF;
rommem[16345] <= 16'hFFFF;
rommem[16346] <= 16'hFFFF;
rommem[16347] <= 16'hFFFF;
rommem[16348] <= 16'hFFFF;
rommem[16349] <= 16'hFFFF;
rommem[16350] <= 16'hFFFF;
rommem[16351] <= 16'hFFFF;
rommem[16352] <= 16'hFFFF;
rommem[16353] <= 16'hFFFF;
rommem[16354] <= 16'hFFFF;
rommem[16355] <= 16'hFFFF;
rommem[16356] <= 16'hFFFF;
rommem[16357] <= 16'hFFFF;
rommem[16358] <= 16'hFFFF;
rommem[16359] <= 16'hFFFF;
rommem[16360] <= 16'hFFFF;
rommem[16361] <= 16'hFFFF;
rommem[16362] <= 16'hFFFF;
rommem[16363] <= 16'hFFFF;
rommem[16364] <= 16'hFFFF;
rommem[16365] <= 16'hFFFF;
rommem[16366] <= 16'hFFFF;
rommem[16367] <= 16'hFFFF;
rommem[16368] <= 16'hFFFF;
rommem[16369] <= 16'hFFFF;
rommem[16370] <= 16'hFFFF;
rommem[16371] <= 16'hFFFF;
rommem[16372] <= 16'hFFFF;
rommem[16373] <= 16'hFFFF;
rommem[16374] <= 16'hFFFF;
rommem[16375] <= 16'hFFFF;
rommem[16376] <= 16'hFFFF;
rommem[16377] <= 16'hFFFF;
rommem[16378] <= 16'hFFFF;
rommem[16379] <= 16'hFFFF;
rommem[16380] <= 16'hFFFF;
rommem[16381] <= 16'hFFFF;
rommem[16382] <= 16'hFFFF;
rommem[16383] <= 16'hFFFF;
rommem[16384] <= 16'hFFFF;
rommem[16385] <= 16'hFFFF;
rommem[16386] <= 16'hFFFF;
rommem[16387] <= 16'hFFFF;
rommem[16388] <= 16'hFFFF;
rommem[16389] <= 16'hFFFF;
rommem[16390] <= 16'hFFFF;
rommem[16391] <= 16'hFFFF;
rommem[16392] <= 16'hFFFF;
rommem[16393] <= 16'hFFFF;
rommem[16394] <= 16'hFFFF;
rommem[16395] <= 16'hFFFF;
rommem[16396] <= 16'hFFFF;
rommem[16397] <= 16'hFFFF;
rommem[16398] <= 16'hFFFF;
rommem[16399] <= 16'hFFFF;
rommem[16400] <= 16'hFFFF;
rommem[16401] <= 16'hFFFF;
rommem[16402] <= 16'hFFFF;
rommem[16403] <= 16'hFFFF;
rommem[16404] <= 16'hFFFF;
rommem[16405] <= 16'hFFFF;
rommem[16406] <= 16'hFFFF;
rommem[16407] <= 16'hFFFF;
rommem[16408] <= 16'hFFFF;
rommem[16409] <= 16'hFFFF;
rommem[16410] <= 16'hFFFF;
rommem[16411] <= 16'hFFFF;
rommem[16412] <= 16'hFFFF;
rommem[16413] <= 16'hFFFF;
rommem[16414] <= 16'hFFFF;
rommem[16415] <= 16'hFFFF;
rommem[16416] <= 16'hFFFF;
rommem[16417] <= 16'hFFFF;
rommem[16418] <= 16'hFFFF;
rommem[16419] <= 16'hFFFF;
rommem[16420] <= 16'hFFFF;
rommem[16421] <= 16'hFFFF;
rommem[16422] <= 16'hFFFF;
rommem[16423] <= 16'hFFFF;
rommem[16424] <= 16'hFFFF;
rommem[16425] <= 16'hFFFF;
rommem[16426] <= 16'hFFFF;
rommem[16427] <= 16'hFFFF;
rommem[16428] <= 16'hFFFF;
rommem[16429] <= 16'hFFFF;
rommem[16430] <= 16'hFFFF;
rommem[16431] <= 16'hFFFF;
rommem[16432] <= 16'hFFFF;
rommem[16433] <= 16'hFFFF;
rommem[16434] <= 16'hFFFF;
rommem[16435] <= 16'hFFFF;
rommem[16436] <= 16'hFFFF;
rommem[16437] <= 16'hFFFF;
rommem[16438] <= 16'hFFFF;
rommem[16439] <= 16'hFFFF;
rommem[16440] <= 16'hFFFF;
rommem[16441] <= 16'hFFFF;
rommem[16442] <= 16'hFFFF;
rommem[16443] <= 16'hFFFF;
rommem[16444] <= 16'hFFFF;
rommem[16445] <= 16'hFFFF;
rommem[16446] <= 16'hFFFF;
rommem[16447] <= 16'hFFFF;
rommem[16448] <= 16'hFFFF;
rommem[16449] <= 16'hFFFF;
rommem[16450] <= 16'hFFFF;
rommem[16451] <= 16'hFFFF;
rommem[16452] <= 16'hFFFF;
rommem[16453] <= 16'hFFFF;
rommem[16454] <= 16'hFFFF;
rommem[16455] <= 16'hFFFF;
rommem[16456] <= 16'hFFFF;
rommem[16457] <= 16'hFFFF;
rommem[16458] <= 16'hFFFF;
rommem[16459] <= 16'hFFFF;
rommem[16460] <= 16'hFFFF;
rommem[16461] <= 16'hFFFF;
rommem[16462] <= 16'hFFFF;
rommem[16463] <= 16'hFFFF;
rommem[16464] <= 16'hFFFF;
rommem[16465] <= 16'hFFFF;
rommem[16466] <= 16'hFFFF;
rommem[16467] <= 16'hFFFF;
rommem[16468] <= 16'hFFFF;
rommem[16469] <= 16'hFFFF;
rommem[16470] <= 16'hFFFF;
rommem[16471] <= 16'hFFFF;
rommem[16472] <= 16'hFFFF;
rommem[16473] <= 16'hFFFF;
rommem[16474] <= 16'hFFFF;
rommem[16475] <= 16'hFFFF;
rommem[16476] <= 16'hFFFF;
rommem[16477] <= 16'hFFFF;
rommem[16478] <= 16'hFFFF;
rommem[16479] <= 16'hFFFF;
rommem[16480] <= 16'hFFFF;
rommem[16481] <= 16'hFFFF;
rommem[16482] <= 16'hFFFF;
rommem[16483] <= 16'hFFFF;
rommem[16484] <= 16'hFFFF;
rommem[16485] <= 16'hFFFF;
rommem[16486] <= 16'hFFFF;
rommem[16487] <= 16'hFFFF;
rommem[16488] <= 16'hFFFF;
rommem[16489] <= 16'hFFFF;
rommem[16490] <= 16'hFFFF;
rommem[16491] <= 16'hFFFF;
rommem[16492] <= 16'hFFFF;
rommem[16493] <= 16'hFFFF;
rommem[16494] <= 16'hFFFF;
rommem[16495] <= 16'hFFFF;
rommem[16496] <= 16'hFFFF;
rommem[16497] <= 16'hFFFF;
rommem[16498] <= 16'hFFFF;
rommem[16499] <= 16'hFFFF;
rommem[16500] <= 16'hFFFF;
rommem[16501] <= 16'hFFFF;
rommem[16502] <= 16'hFFFF;
rommem[16503] <= 16'hFFFF;
rommem[16504] <= 16'hFFFF;
rommem[16505] <= 16'hFFFF;
rommem[16506] <= 16'hFFFF;
rommem[16507] <= 16'hFFFF;
rommem[16508] <= 16'hFFFF;
rommem[16509] <= 16'hFFFF;
rommem[16510] <= 16'hFFFF;
rommem[16511] <= 16'hFFFF;
rommem[16512] <= 16'hFFFF;
rommem[16513] <= 16'hFFFF;
rommem[16514] <= 16'hFFFF;
rommem[16515] <= 16'hFFFF;
rommem[16516] <= 16'hFFFF;
rommem[16517] <= 16'hFFFF;
rommem[16518] <= 16'hFFFF;
rommem[16519] <= 16'hFFFF;
rommem[16520] <= 16'hFFFF;
rommem[16521] <= 16'hFFFF;
rommem[16522] <= 16'hFFFF;
rommem[16523] <= 16'hFFFF;
rommem[16524] <= 16'hFFFF;
rommem[16525] <= 16'hFFFF;
rommem[16526] <= 16'hFFFF;
rommem[16527] <= 16'hFFFF;
rommem[16528] <= 16'hFFFF;
rommem[16529] <= 16'hFFFF;
rommem[16530] <= 16'hFFFF;
rommem[16531] <= 16'hFFFF;
rommem[16532] <= 16'hFFFF;
rommem[16533] <= 16'hFFFF;
rommem[16534] <= 16'hFFFF;
rommem[16535] <= 16'hFFFF;
rommem[16536] <= 16'hFFFF;
rommem[16537] <= 16'hFFFF;
rommem[16538] <= 16'hFFFF;
rommem[16539] <= 16'hFFFF;
rommem[16540] <= 16'hFFFF;
rommem[16541] <= 16'hFFFF;
rommem[16542] <= 16'hFFFF;
rommem[16543] <= 16'hFFFF;
rommem[16544] <= 16'hFFFF;
rommem[16545] <= 16'hFFFF;
rommem[16546] <= 16'hFFFF;
rommem[16547] <= 16'hFFFF;
rommem[16548] <= 16'hFFFF;
rommem[16549] <= 16'hFFFF;
rommem[16550] <= 16'hFFFF;
rommem[16551] <= 16'hFFFF;
rommem[16552] <= 16'hFFFF;
rommem[16553] <= 16'hFFFF;
rommem[16554] <= 16'hFFFF;
rommem[16555] <= 16'hFFFF;
rommem[16556] <= 16'hFFFF;
rommem[16557] <= 16'hFFFF;
rommem[16558] <= 16'hFFFF;
rommem[16559] <= 16'hFFFF;
rommem[16560] <= 16'hFFFF;
rommem[16561] <= 16'hFFFF;
rommem[16562] <= 16'hFFFF;
rommem[16563] <= 16'hFFFF;
rommem[16564] <= 16'hFFFF;
rommem[16565] <= 16'hFFFF;
rommem[16566] <= 16'hFFFF;
rommem[16567] <= 16'hFFFF;
rommem[16568] <= 16'hFFFF;
rommem[16569] <= 16'hFFFF;
rommem[16570] <= 16'hFFFF;
rommem[16571] <= 16'hFFFF;
rommem[16572] <= 16'hFFFF;
rommem[16573] <= 16'hFFFF;
rommem[16574] <= 16'hFFFF;
rommem[16575] <= 16'hFFFF;
rommem[16576] <= 16'hFFFF;
rommem[16577] <= 16'hFFFF;
rommem[16578] <= 16'hFFFF;
rommem[16579] <= 16'hFFFF;
rommem[16580] <= 16'hFFFF;
rommem[16581] <= 16'hFFFF;
rommem[16582] <= 16'hFFFF;
rommem[16583] <= 16'hFFFF;
rommem[16584] <= 16'hFFFF;
rommem[16585] <= 16'hFFFF;
rommem[16586] <= 16'hFFFF;
rommem[16587] <= 16'hFFFF;
rommem[16588] <= 16'hFFFF;
rommem[16589] <= 16'hFFFF;
rommem[16590] <= 16'hFFFF;
rommem[16591] <= 16'hFFFF;
rommem[16592] <= 16'hFFFF;
rommem[16593] <= 16'hFFFF;
rommem[16594] <= 16'hFFFF;
rommem[16595] <= 16'hFFFF;
rommem[16596] <= 16'hFFFF;
rommem[16597] <= 16'hFFFF;
rommem[16598] <= 16'hFFFF;
rommem[16599] <= 16'hFFFF;
rommem[16600] <= 16'hFFFF;
rommem[16601] <= 16'hFFFF;
rommem[16602] <= 16'hFFFF;
rommem[16603] <= 16'hFFFF;
rommem[16604] <= 16'hFFFF;
rommem[16605] <= 16'hFFFF;
rommem[16606] <= 16'hFFFF;
rommem[16607] <= 16'hFFFF;
rommem[16608] <= 16'hFFFF;
rommem[16609] <= 16'hFFFF;
rommem[16610] <= 16'hFFFF;
rommem[16611] <= 16'hFFFF;
rommem[16612] <= 16'hFFFF;
rommem[16613] <= 16'hFFFF;
rommem[16614] <= 16'hFFFF;
rommem[16615] <= 16'hFFFF;
rommem[16616] <= 16'hFFFF;
rommem[16617] <= 16'hFFFF;
rommem[16618] <= 16'hFFFF;
rommem[16619] <= 16'hFFFF;
rommem[16620] <= 16'hFFFF;
rommem[16621] <= 16'hFFFF;
rommem[16622] <= 16'hFFFF;
rommem[16623] <= 16'hFFFF;
rommem[16624] <= 16'hFFFF;
rommem[16625] <= 16'hFFFF;
rommem[16626] <= 16'hFFFF;
rommem[16627] <= 16'hFFFF;
rommem[16628] <= 16'hFFFF;
rommem[16629] <= 16'hFFFF;
rommem[16630] <= 16'hFFFF;
rommem[16631] <= 16'hFFFF;
rommem[16632] <= 16'hFFFF;
rommem[16633] <= 16'hFFFF;
rommem[16634] <= 16'hFFFF;
rommem[16635] <= 16'hFFFF;
rommem[16636] <= 16'hFFFF;
rommem[16637] <= 16'hFFFF;
rommem[16638] <= 16'hFFFF;
rommem[16639] <= 16'hFFFF;
rommem[16640] <= 16'hFFFF;
rommem[16641] <= 16'hFFFF;
rommem[16642] <= 16'hFFFF;
rommem[16643] <= 16'hFFFF;
rommem[16644] <= 16'hFFFF;
rommem[16645] <= 16'hFFFF;
rommem[16646] <= 16'hFFFF;
rommem[16647] <= 16'hFFFF;
rommem[16648] <= 16'hFFFF;
rommem[16649] <= 16'hFFFF;
rommem[16650] <= 16'hFFFF;
rommem[16651] <= 16'hFFFF;
rommem[16652] <= 16'hFFFF;
rommem[16653] <= 16'hFFFF;
rommem[16654] <= 16'hFFFF;
rommem[16655] <= 16'hFFFF;
rommem[16656] <= 16'hFFFF;
rommem[16657] <= 16'hFFFF;
rommem[16658] <= 16'hFFFF;
rommem[16659] <= 16'hFFFF;
rommem[16660] <= 16'hFFFF;
rommem[16661] <= 16'hFFFF;
rommem[16662] <= 16'hFFFF;
rommem[16663] <= 16'hFFFF;
rommem[16664] <= 16'hFFFF;
rommem[16665] <= 16'hFFFF;
rommem[16666] <= 16'hFFFF;
rommem[16667] <= 16'hFFFF;
rommem[16668] <= 16'hFFFF;
rommem[16669] <= 16'hFFFF;
rommem[16670] <= 16'hFFFF;
rommem[16671] <= 16'hFFFF;
rommem[16672] <= 16'hFFFF;
rommem[16673] <= 16'hFFFF;
rommem[16674] <= 16'hFFFF;
rommem[16675] <= 16'hFFFF;
rommem[16676] <= 16'hFFFF;
rommem[16677] <= 16'hFFFF;
rommem[16678] <= 16'hFFFF;
rommem[16679] <= 16'hFFFF;
rommem[16680] <= 16'hFFFF;
rommem[16681] <= 16'hFFFF;
rommem[16682] <= 16'hFFFF;
rommem[16683] <= 16'hFFFF;
rommem[16684] <= 16'hFFFF;
rommem[16685] <= 16'hFFFF;
rommem[16686] <= 16'hFFFF;
rommem[16687] <= 16'hFFFF;
rommem[16688] <= 16'hFFFF;
rommem[16689] <= 16'hFFFF;
rommem[16690] <= 16'hFFFF;
rommem[16691] <= 16'hFFFF;
rommem[16692] <= 16'hFFFF;
rommem[16693] <= 16'hFFFF;
rommem[16694] <= 16'hFFFF;
rommem[16695] <= 16'hFFFF;
rommem[16696] <= 16'hFFFF;
rommem[16697] <= 16'hFFFF;
rommem[16698] <= 16'hFFFF;
rommem[16699] <= 16'hFFFF;
rommem[16700] <= 16'hFFFF;
rommem[16701] <= 16'hFFFF;
rommem[16702] <= 16'hFFFF;
rommem[16703] <= 16'hFFFF;
rommem[16704] <= 16'hFFFF;
rommem[16705] <= 16'hFFFF;
rommem[16706] <= 16'hFFFF;
rommem[16707] <= 16'hFFFF;
rommem[16708] <= 16'hFFFF;
rommem[16709] <= 16'hFFFF;
rommem[16710] <= 16'hFFFF;
rommem[16711] <= 16'hFFFF;
rommem[16712] <= 16'hFFFF;
rommem[16713] <= 16'hFFFF;
rommem[16714] <= 16'hFFFF;
rommem[16715] <= 16'hFFFF;
rommem[16716] <= 16'hFFFF;
rommem[16717] <= 16'hFFFF;
rommem[16718] <= 16'hFFFF;
rommem[16719] <= 16'hFFFF;
rommem[16720] <= 16'hFFFF;
rommem[16721] <= 16'hFFFF;
rommem[16722] <= 16'hFFFF;
rommem[16723] <= 16'hFFFF;
rommem[16724] <= 16'hFFFF;
rommem[16725] <= 16'hFFFF;
rommem[16726] <= 16'hFFFF;
rommem[16727] <= 16'hFFFF;
rommem[16728] <= 16'hFFFF;
rommem[16729] <= 16'hFFFF;
rommem[16730] <= 16'hFFFF;
rommem[16731] <= 16'hFFFF;
rommem[16732] <= 16'hFFFF;
rommem[16733] <= 16'hFFFF;
rommem[16734] <= 16'hFFFF;
rommem[16735] <= 16'hFFFF;
rommem[16736] <= 16'hFFFF;
rommem[16737] <= 16'hFFFF;
rommem[16738] <= 16'hFFFF;
rommem[16739] <= 16'hFFFF;
rommem[16740] <= 16'hFFFF;
rommem[16741] <= 16'hFFFF;
rommem[16742] <= 16'hFFFF;
rommem[16743] <= 16'hFFFF;
rommem[16744] <= 16'hFFFF;
rommem[16745] <= 16'hFFFF;
rommem[16746] <= 16'hFFFF;
rommem[16747] <= 16'hFFFF;
rommem[16748] <= 16'hFFFF;
rommem[16749] <= 16'hFFFF;
rommem[16750] <= 16'hFFFF;
rommem[16751] <= 16'hFFFF;
rommem[16752] <= 16'hFFFF;
rommem[16753] <= 16'hFFFF;
rommem[16754] <= 16'hFFFF;
rommem[16755] <= 16'hFFFF;
rommem[16756] <= 16'hFFFF;
rommem[16757] <= 16'hFFFF;
rommem[16758] <= 16'hFFFF;
rommem[16759] <= 16'hFFFF;
rommem[16760] <= 16'hFFFF;
rommem[16761] <= 16'hFFFF;
rommem[16762] <= 16'hFFFF;
rommem[16763] <= 16'hFFFF;
rommem[16764] <= 16'hFFFF;
rommem[16765] <= 16'hFFFF;
rommem[16766] <= 16'hFFFF;
rommem[16767] <= 16'hFFFF;
rommem[16768] <= 16'hFFFF;
rommem[16769] <= 16'hFFFF;
rommem[16770] <= 16'hFFFF;
rommem[16771] <= 16'hFFFF;
rommem[16772] <= 16'hFFFF;
rommem[16773] <= 16'hFFFF;
rommem[16774] <= 16'hFFFF;
rommem[16775] <= 16'hFFFF;
rommem[16776] <= 16'hFFFF;
rommem[16777] <= 16'hFFFF;
rommem[16778] <= 16'hFFFF;
rommem[16779] <= 16'hFFFF;
rommem[16780] <= 16'hFFFF;
rommem[16781] <= 16'hFFFF;
rommem[16782] <= 16'hFFFF;
rommem[16783] <= 16'hFFFF;
rommem[16784] <= 16'hFFFF;
rommem[16785] <= 16'hFFFF;
rommem[16786] <= 16'hFFFF;
rommem[16787] <= 16'hFFFF;
rommem[16788] <= 16'hFFFF;
rommem[16789] <= 16'hFFFF;
rommem[16790] <= 16'hFFFF;
rommem[16791] <= 16'hFFFF;
rommem[16792] <= 16'hFFFF;
rommem[16793] <= 16'hFFFF;
rommem[16794] <= 16'hFFFF;
rommem[16795] <= 16'hFFFF;
rommem[16796] <= 16'hFFFF;
rommem[16797] <= 16'hFFFF;
rommem[16798] <= 16'hFFFF;
rommem[16799] <= 16'hFFFF;
rommem[16800] <= 16'hFFFF;
rommem[16801] <= 16'hFFFF;
rommem[16802] <= 16'hFFFF;
rommem[16803] <= 16'hFFFF;
rommem[16804] <= 16'hFFFF;
rommem[16805] <= 16'hFFFF;
rommem[16806] <= 16'hFFFF;
rommem[16807] <= 16'hFFFF;
rommem[16808] <= 16'hFFFF;
rommem[16809] <= 16'hFFFF;
rommem[16810] <= 16'hFFFF;
rommem[16811] <= 16'hFFFF;
rommem[16812] <= 16'hFFFF;
rommem[16813] <= 16'hFFFF;
rommem[16814] <= 16'hFFFF;
rommem[16815] <= 16'hFFFF;
rommem[16816] <= 16'hFFFF;
rommem[16817] <= 16'hFFFF;
rommem[16818] <= 16'hFFFF;
rommem[16819] <= 16'hFFFF;
rommem[16820] <= 16'hFFFF;
rommem[16821] <= 16'hFFFF;
rommem[16822] <= 16'hFFFF;
rommem[16823] <= 16'hFFFF;
rommem[16824] <= 16'hFFFF;
rommem[16825] <= 16'hFFFF;
rommem[16826] <= 16'hFFFF;
rommem[16827] <= 16'hFFFF;
rommem[16828] <= 16'hFFFF;
rommem[16829] <= 16'hFFFF;
rommem[16830] <= 16'hFFFF;
rommem[16831] <= 16'hFFFF;
rommem[16832] <= 16'hFFFF;
rommem[16833] <= 16'hFFFF;
rommem[16834] <= 16'hFFFF;
rommem[16835] <= 16'hFFFF;
rommem[16836] <= 16'hFFFF;
rommem[16837] <= 16'hFFFF;
rommem[16838] <= 16'hFFFF;
rommem[16839] <= 16'hFFFF;
rommem[16840] <= 16'hFFFF;
rommem[16841] <= 16'hFFFF;
rommem[16842] <= 16'hFFFF;
rommem[16843] <= 16'hFFFF;
rommem[16844] <= 16'hFFFF;
rommem[16845] <= 16'hFFFF;
rommem[16846] <= 16'hFFFF;
rommem[16847] <= 16'hFFFF;
rommem[16848] <= 16'hFFFF;
rommem[16849] <= 16'hFFFF;
rommem[16850] <= 16'hFFFF;
rommem[16851] <= 16'hFFFF;
rommem[16852] <= 16'hFFFF;
rommem[16853] <= 16'hFFFF;
rommem[16854] <= 16'hFFFF;
rommem[16855] <= 16'hFFFF;
rommem[16856] <= 16'hFFFF;
rommem[16857] <= 16'hFFFF;
rommem[16858] <= 16'hFFFF;
rommem[16859] <= 16'hFFFF;
rommem[16860] <= 16'hFFFF;
rommem[16861] <= 16'hFFFF;
rommem[16862] <= 16'hFFFF;
rommem[16863] <= 16'hFFFF;
rommem[16864] <= 16'hFFFF;
rommem[16865] <= 16'hFFFF;
rommem[16866] <= 16'hFFFF;
rommem[16867] <= 16'hFFFF;
rommem[16868] <= 16'hFFFF;
rommem[16869] <= 16'hFFFF;
rommem[16870] <= 16'hFFFF;
rommem[16871] <= 16'hFFFF;
rommem[16872] <= 16'hFFFF;
rommem[16873] <= 16'hFFFF;
rommem[16874] <= 16'hFFFF;
rommem[16875] <= 16'hFFFF;
rommem[16876] <= 16'hFFFF;
rommem[16877] <= 16'hFFFF;
rommem[16878] <= 16'hFFFF;
rommem[16879] <= 16'hFFFF;
rommem[16880] <= 16'hFFFF;
rommem[16881] <= 16'hFFFF;
rommem[16882] <= 16'hFFFF;
rommem[16883] <= 16'hFFFF;
rommem[16884] <= 16'hFFFF;
rommem[16885] <= 16'hFFFF;
rommem[16886] <= 16'hFFFF;
rommem[16887] <= 16'hFFFF;
rommem[16888] <= 16'hFFFF;
rommem[16889] <= 16'hFFFF;
rommem[16890] <= 16'hFFFF;
rommem[16891] <= 16'hFFFF;
rommem[16892] <= 16'hFFFF;
rommem[16893] <= 16'hFFFF;
rommem[16894] <= 16'hFFFF;
rommem[16895] <= 16'hFFFF;
rommem[16896] <= 16'hFFFF;
rommem[16897] <= 16'hFFFF;
rommem[16898] <= 16'hFFFF;
rommem[16899] <= 16'hFFFF;
rommem[16900] <= 16'hFFFF;
rommem[16901] <= 16'hFFFF;
rommem[16902] <= 16'hFFFF;
rommem[16903] <= 16'hFFFF;
rommem[16904] <= 16'hFFFF;
rommem[16905] <= 16'hFFFF;
rommem[16906] <= 16'hFFFF;
rommem[16907] <= 16'hFFFF;
rommem[16908] <= 16'hFFFF;
rommem[16909] <= 16'hFFFF;
rommem[16910] <= 16'hFFFF;
rommem[16911] <= 16'hFFFF;
rommem[16912] <= 16'hFFFF;
rommem[16913] <= 16'hFFFF;
rommem[16914] <= 16'hFFFF;
rommem[16915] <= 16'hFFFF;
rommem[16916] <= 16'hFFFF;
rommem[16917] <= 16'hFFFF;
rommem[16918] <= 16'hFFFF;
rommem[16919] <= 16'hFFFF;
rommem[16920] <= 16'hFFFF;
rommem[16921] <= 16'hFFFF;
rommem[16922] <= 16'hFFFF;
rommem[16923] <= 16'hFFFF;
rommem[16924] <= 16'hFFFF;
rommem[16925] <= 16'hFFFF;
rommem[16926] <= 16'hFFFF;
rommem[16927] <= 16'hFFFF;
rommem[16928] <= 16'hFFFF;
rommem[16929] <= 16'hFFFF;
rommem[16930] <= 16'hFFFF;
rommem[16931] <= 16'hFFFF;
rommem[16932] <= 16'hFFFF;
rommem[16933] <= 16'hFFFF;
rommem[16934] <= 16'hFFFF;
rommem[16935] <= 16'hFFFF;
rommem[16936] <= 16'hFFFF;
rommem[16937] <= 16'hFFFF;
rommem[16938] <= 16'hFFFF;
rommem[16939] <= 16'hFFFF;
rommem[16940] <= 16'hFFFF;
rommem[16941] <= 16'hFFFF;
rommem[16942] <= 16'hFFFF;
rommem[16943] <= 16'hFFFF;
rommem[16944] <= 16'hFFFF;
rommem[16945] <= 16'hFFFF;
rommem[16946] <= 16'hFFFF;
rommem[16947] <= 16'hFFFF;
rommem[16948] <= 16'hFFFF;
rommem[16949] <= 16'hFFFF;
rommem[16950] <= 16'hFFFF;
rommem[16951] <= 16'hFFFF;
rommem[16952] <= 16'hFFFF;
rommem[16953] <= 16'hFFFF;
rommem[16954] <= 16'hFFFF;
rommem[16955] <= 16'hFFFF;
rommem[16956] <= 16'hFFFF;
rommem[16957] <= 16'hFFFF;
rommem[16958] <= 16'hFFFF;
rommem[16959] <= 16'hFFFF;
rommem[16960] <= 16'hFFFF;
rommem[16961] <= 16'hFFFF;
rommem[16962] <= 16'hFFFF;
rommem[16963] <= 16'hFFFF;
rommem[16964] <= 16'hFFFF;
rommem[16965] <= 16'hFFFF;
rommem[16966] <= 16'hFFFF;
rommem[16967] <= 16'hFFFF;
rommem[16968] <= 16'hFFFF;
rommem[16969] <= 16'hFFFF;
rommem[16970] <= 16'hFFFF;
rommem[16971] <= 16'hFFFF;
rommem[16972] <= 16'hFFFF;
rommem[16973] <= 16'hFFFF;
rommem[16974] <= 16'hFFFF;
rommem[16975] <= 16'hFFFF;
rommem[16976] <= 16'hFFFF;
rommem[16977] <= 16'hFFFF;
rommem[16978] <= 16'hFFFF;
rommem[16979] <= 16'hFFFF;
rommem[16980] <= 16'hFFFF;
rommem[16981] <= 16'hFFFF;
rommem[16982] <= 16'hFFFF;
rommem[16983] <= 16'hFFFF;
rommem[16984] <= 16'hFFFF;
rommem[16985] <= 16'hFFFF;
rommem[16986] <= 16'hFFFF;
rommem[16987] <= 16'hFFFF;
rommem[16988] <= 16'hFFFF;
rommem[16989] <= 16'hFFFF;
rommem[16990] <= 16'hFFFF;
rommem[16991] <= 16'hFFFF;
rommem[16992] <= 16'hFFFF;
rommem[16993] <= 16'hFFFF;
rommem[16994] <= 16'hFFFF;
rommem[16995] <= 16'hFFFF;
rommem[16996] <= 16'hFFFF;
rommem[16997] <= 16'hFFFF;
rommem[16998] <= 16'hFFFF;
rommem[16999] <= 16'hFFFF;
rommem[17000] <= 16'hFFFF;
rommem[17001] <= 16'hFFFF;
rommem[17002] <= 16'hFFFF;
rommem[17003] <= 16'hFFFF;
rommem[17004] <= 16'hFFFF;
rommem[17005] <= 16'hFFFF;
rommem[17006] <= 16'hFFFF;
rommem[17007] <= 16'hFFFF;
rommem[17008] <= 16'hFFFF;
rommem[17009] <= 16'hFFFF;
rommem[17010] <= 16'hFFFF;
rommem[17011] <= 16'hFFFF;
rommem[17012] <= 16'hFFFF;
rommem[17013] <= 16'hFFFF;
rommem[17014] <= 16'hFFFF;
rommem[17015] <= 16'hFFFF;
rommem[17016] <= 16'hFFFF;
rommem[17017] <= 16'hFFFF;
rommem[17018] <= 16'hFFFF;
rommem[17019] <= 16'hFFFF;
rommem[17020] <= 16'hFFFF;
rommem[17021] <= 16'hFFFF;
rommem[17022] <= 16'hFFFF;
rommem[17023] <= 16'hFFFF;
rommem[17024] <= 16'hFFFF;
rommem[17025] <= 16'hFFFF;
rommem[17026] <= 16'hFFFF;
rommem[17027] <= 16'hFFFF;
rommem[17028] <= 16'hFFFF;
rommem[17029] <= 16'hFFFF;
rommem[17030] <= 16'hFFFF;
rommem[17031] <= 16'hFFFF;
rommem[17032] <= 16'hFFFF;
rommem[17033] <= 16'hFFFF;
rommem[17034] <= 16'hFFFF;
rommem[17035] <= 16'hFFFF;
rommem[17036] <= 16'hFFFF;
rommem[17037] <= 16'hFFFF;
rommem[17038] <= 16'hFFFF;
rommem[17039] <= 16'hFFFF;
rommem[17040] <= 16'hFFFF;
rommem[17041] <= 16'hFFFF;
rommem[17042] <= 16'hFFFF;
rommem[17043] <= 16'hFFFF;
rommem[17044] <= 16'hFFFF;
rommem[17045] <= 16'hFFFF;
rommem[17046] <= 16'hFFFF;
rommem[17047] <= 16'hFFFF;
rommem[17048] <= 16'hFFFF;
rommem[17049] <= 16'hFFFF;
rommem[17050] <= 16'hFFFF;
rommem[17051] <= 16'hFFFF;
rommem[17052] <= 16'hFFFF;
rommem[17053] <= 16'hFFFF;
rommem[17054] <= 16'hFFFF;
rommem[17055] <= 16'hFFFF;
rommem[17056] <= 16'hFFFF;
rommem[17057] <= 16'hFFFF;
rommem[17058] <= 16'hFFFF;
rommem[17059] <= 16'hFFFF;
rommem[17060] <= 16'hFFFF;
rommem[17061] <= 16'hFFFF;
rommem[17062] <= 16'hFFFF;
rommem[17063] <= 16'hFFFF;
rommem[17064] <= 16'hFFFF;
rommem[17065] <= 16'hFFFF;
rommem[17066] <= 16'hFFFF;
rommem[17067] <= 16'hFFFF;
rommem[17068] <= 16'hFFFF;
rommem[17069] <= 16'hFFFF;
rommem[17070] <= 16'hFFFF;
rommem[17071] <= 16'hFFFF;
rommem[17072] <= 16'hFFFF;
rommem[17073] <= 16'hFFFF;
rommem[17074] <= 16'hFFFF;
rommem[17075] <= 16'hFFFF;
rommem[17076] <= 16'hFFFF;
rommem[17077] <= 16'hFFFF;
rommem[17078] <= 16'hFFFF;
rommem[17079] <= 16'hFFFF;
rommem[17080] <= 16'hFFFF;
rommem[17081] <= 16'hFFFF;
rommem[17082] <= 16'hFFFF;
rommem[17083] <= 16'hFFFF;
rommem[17084] <= 16'hFFFF;
rommem[17085] <= 16'hFFFF;
rommem[17086] <= 16'hFFFF;
rommem[17087] <= 16'hFFFF;
rommem[17088] <= 16'hFFFF;
rommem[17089] <= 16'hFFFF;
rommem[17090] <= 16'hFFFF;
rommem[17091] <= 16'hFFFF;
rommem[17092] <= 16'hFFFF;
rommem[17093] <= 16'hFFFF;
rommem[17094] <= 16'hFFFF;
rommem[17095] <= 16'hFFFF;
rommem[17096] <= 16'hFFFF;
rommem[17097] <= 16'hFFFF;
rommem[17098] <= 16'hFFFF;
rommem[17099] <= 16'hFFFF;
rommem[17100] <= 16'hFFFF;
rommem[17101] <= 16'hFFFF;
rommem[17102] <= 16'hFFFF;
rommem[17103] <= 16'hFFFF;
rommem[17104] <= 16'hFFFF;
rommem[17105] <= 16'hFFFF;
rommem[17106] <= 16'hFFFF;
rommem[17107] <= 16'hFFFF;
rommem[17108] <= 16'hFFFF;
rommem[17109] <= 16'hFFFF;
rommem[17110] <= 16'hFFFF;
rommem[17111] <= 16'hFFFF;
rommem[17112] <= 16'hFFFF;
rommem[17113] <= 16'hFFFF;
rommem[17114] <= 16'hFFFF;
rommem[17115] <= 16'hFFFF;
rommem[17116] <= 16'hFFFF;
rommem[17117] <= 16'hFFFF;
rommem[17118] <= 16'hFFFF;
rommem[17119] <= 16'hFFFF;
rommem[17120] <= 16'hFFFF;
rommem[17121] <= 16'hFFFF;
rommem[17122] <= 16'hFFFF;
rommem[17123] <= 16'hFFFF;
rommem[17124] <= 16'hFFFF;
rommem[17125] <= 16'hFFFF;
rommem[17126] <= 16'hFFFF;
rommem[17127] <= 16'hFFFF;
rommem[17128] <= 16'hFFFF;
rommem[17129] <= 16'hFFFF;
rommem[17130] <= 16'hFFFF;
rommem[17131] <= 16'hFFFF;
rommem[17132] <= 16'hFFFF;
rommem[17133] <= 16'hFFFF;
rommem[17134] <= 16'hFFFF;
rommem[17135] <= 16'hFFFF;
rommem[17136] <= 16'hFFFF;
rommem[17137] <= 16'hFFFF;
rommem[17138] <= 16'hFFFF;
rommem[17139] <= 16'hFFFF;
rommem[17140] <= 16'hFFFF;
rommem[17141] <= 16'hFFFF;
rommem[17142] <= 16'hFFFF;
rommem[17143] <= 16'hFFFF;
rommem[17144] <= 16'hFFFF;
rommem[17145] <= 16'hFFFF;
rommem[17146] <= 16'hFFFF;
rommem[17147] <= 16'hFFFF;
rommem[17148] <= 16'hFFFF;
rommem[17149] <= 16'hFFFF;
rommem[17150] <= 16'hFFFF;
rommem[17151] <= 16'hFFFF;
rommem[17152] <= 16'hFFFF;
rommem[17153] <= 16'hFFFF;
rommem[17154] <= 16'hFFFF;
rommem[17155] <= 16'hFFFF;
rommem[17156] <= 16'hFFFF;
rommem[17157] <= 16'hFFFF;
rommem[17158] <= 16'hFFFF;
rommem[17159] <= 16'hFFFF;
rommem[17160] <= 16'hFFFF;
rommem[17161] <= 16'hFFFF;
rommem[17162] <= 16'hFFFF;
rommem[17163] <= 16'hFFFF;
rommem[17164] <= 16'hFFFF;
rommem[17165] <= 16'hFFFF;
rommem[17166] <= 16'hFFFF;
rommem[17167] <= 16'hFFFF;
rommem[17168] <= 16'hFFFF;
rommem[17169] <= 16'hFFFF;
rommem[17170] <= 16'hFFFF;
rommem[17171] <= 16'hFFFF;
rommem[17172] <= 16'hFFFF;
rommem[17173] <= 16'hFFFF;
rommem[17174] <= 16'hFFFF;
rommem[17175] <= 16'hFFFF;
rommem[17176] <= 16'hFFFF;
rommem[17177] <= 16'hFFFF;
rommem[17178] <= 16'hFFFF;
rommem[17179] <= 16'hFFFF;
rommem[17180] <= 16'hFFFF;
rommem[17181] <= 16'hFFFF;
rommem[17182] <= 16'hFFFF;
rommem[17183] <= 16'hFFFF;
rommem[17184] <= 16'hFFFF;
rommem[17185] <= 16'hFFFF;
rommem[17186] <= 16'hFFFF;
rommem[17187] <= 16'hFFFF;
rommem[17188] <= 16'hFFFF;
rommem[17189] <= 16'hFFFF;
rommem[17190] <= 16'hFFFF;
rommem[17191] <= 16'hFFFF;
rommem[17192] <= 16'hFFFF;
rommem[17193] <= 16'hFFFF;
rommem[17194] <= 16'hFFFF;
rommem[17195] <= 16'hFFFF;
rommem[17196] <= 16'hFFFF;
rommem[17197] <= 16'hFFFF;
rommem[17198] <= 16'hFFFF;
rommem[17199] <= 16'hFFFF;
rommem[17200] <= 16'hFFFF;
rommem[17201] <= 16'hFFFF;
rommem[17202] <= 16'hFFFF;
rommem[17203] <= 16'hFFFF;
rommem[17204] <= 16'hFFFF;
rommem[17205] <= 16'hFFFF;
rommem[17206] <= 16'hFFFF;
rommem[17207] <= 16'hFFFF;
rommem[17208] <= 16'hFFFF;
rommem[17209] <= 16'hFFFF;
rommem[17210] <= 16'hFFFF;
rommem[17211] <= 16'hFFFF;
rommem[17212] <= 16'hFFFF;
rommem[17213] <= 16'hFFFF;
rommem[17214] <= 16'hFFFF;
rommem[17215] <= 16'hFFFF;
rommem[17216] <= 16'hFFFF;
rommem[17217] <= 16'hFFFF;
rommem[17218] <= 16'hFFFF;
rommem[17219] <= 16'hFFFF;
rommem[17220] <= 16'hFFFF;
rommem[17221] <= 16'hFFFF;
rommem[17222] <= 16'hFFFF;
rommem[17223] <= 16'hFFFF;
rommem[17224] <= 16'hFFFF;
rommem[17225] <= 16'hFFFF;
rommem[17226] <= 16'hFFFF;
rommem[17227] <= 16'hFFFF;
rommem[17228] <= 16'hFFFF;
rommem[17229] <= 16'hFFFF;
rommem[17230] <= 16'hFFFF;
rommem[17231] <= 16'hFFFF;
rommem[17232] <= 16'hFFFF;
rommem[17233] <= 16'hFFFF;
rommem[17234] <= 16'hFFFF;
rommem[17235] <= 16'hFFFF;
rommem[17236] <= 16'hFFFF;
rommem[17237] <= 16'hFFFF;
rommem[17238] <= 16'hFFFF;
rommem[17239] <= 16'hFFFF;
rommem[17240] <= 16'hFFFF;
rommem[17241] <= 16'hFFFF;
rommem[17242] <= 16'hFFFF;
rommem[17243] <= 16'hFFFF;
rommem[17244] <= 16'hFFFF;
rommem[17245] <= 16'hFFFF;
rommem[17246] <= 16'hFFFF;
rommem[17247] <= 16'hFFFF;
rommem[17248] <= 16'hFFFF;
rommem[17249] <= 16'hFFFF;
rommem[17250] <= 16'hFFFF;
rommem[17251] <= 16'hFFFF;
rommem[17252] <= 16'hFFFF;
rommem[17253] <= 16'hFFFF;
rommem[17254] <= 16'hFFFF;
rommem[17255] <= 16'hFFFF;
rommem[17256] <= 16'hFFFF;
rommem[17257] <= 16'hFFFF;
rommem[17258] <= 16'hFFFF;
rommem[17259] <= 16'hFFFF;
rommem[17260] <= 16'hFFFF;
rommem[17261] <= 16'hFFFF;
rommem[17262] <= 16'hFFFF;
rommem[17263] <= 16'hFFFF;
rommem[17264] <= 16'hFFFF;
rommem[17265] <= 16'hFFFF;
rommem[17266] <= 16'hFFFF;
rommem[17267] <= 16'hFFFF;
rommem[17268] <= 16'hFFFF;
rommem[17269] <= 16'hFFFF;
rommem[17270] <= 16'hFFFF;
rommem[17271] <= 16'hFFFF;
rommem[17272] <= 16'hFFFF;
rommem[17273] <= 16'hFFFF;
rommem[17274] <= 16'hFFFF;
rommem[17275] <= 16'hFFFF;
rommem[17276] <= 16'hFFFF;
rommem[17277] <= 16'hFFFF;
rommem[17278] <= 16'hFFFF;
rommem[17279] <= 16'hFFFF;
rommem[17280] <= 16'hFFFF;
rommem[17281] <= 16'hFFFF;
rommem[17282] <= 16'hFFFF;
rommem[17283] <= 16'hFFFF;
rommem[17284] <= 16'hFFFF;
rommem[17285] <= 16'hFFFF;
rommem[17286] <= 16'hFFFF;
rommem[17287] <= 16'hFFFF;
rommem[17288] <= 16'hFFFF;
rommem[17289] <= 16'hFFFF;
rommem[17290] <= 16'hFFFF;
rommem[17291] <= 16'hFFFF;
rommem[17292] <= 16'hFFFF;
rommem[17293] <= 16'hFFFF;
rommem[17294] <= 16'hFFFF;
rommem[17295] <= 16'hFFFF;
rommem[17296] <= 16'hFFFF;
rommem[17297] <= 16'hFFFF;
rommem[17298] <= 16'hFFFF;
rommem[17299] <= 16'hFFFF;
rommem[17300] <= 16'hFFFF;
rommem[17301] <= 16'hFFFF;
rommem[17302] <= 16'hFFFF;
rommem[17303] <= 16'hFFFF;
rommem[17304] <= 16'hFFFF;
rommem[17305] <= 16'hFFFF;
rommem[17306] <= 16'hFFFF;
rommem[17307] <= 16'hFFFF;
rommem[17308] <= 16'hFFFF;
rommem[17309] <= 16'hFFFF;
rommem[17310] <= 16'hFFFF;
rommem[17311] <= 16'hFFFF;
rommem[17312] <= 16'hFFFF;
rommem[17313] <= 16'hFFFF;
rommem[17314] <= 16'hFFFF;
rommem[17315] <= 16'hFFFF;
rommem[17316] <= 16'hFFFF;
rommem[17317] <= 16'hFFFF;
rommem[17318] <= 16'hFFFF;
rommem[17319] <= 16'hFFFF;
rommem[17320] <= 16'hFFFF;
rommem[17321] <= 16'hFFFF;
rommem[17322] <= 16'hFFFF;
rommem[17323] <= 16'hFFFF;
rommem[17324] <= 16'hFFFF;
rommem[17325] <= 16'hFFFF;
rommem[17326] <= 16'hFFFF;
rommem[17327] <= 16'hFFFF;
rommem[17328] <= 16'hFFFF;
rommem[17329] <= 16'hFFFF;
rommem[17330] <= 16'hFFFF;
rommem[17331] <= 16'hFFFF;
rommem[17332] <= 16'hFFFF;
rommem[17333] <= 16'hFFFF;
rommem[17334] <= 16'hFFFF;
rommem[17335] <= 16'hFFFF;
rommem[17336] <= 16'hFFFF;
rommem[17337] <= 16'hFFFF;
rommem[17338] <= 16'hFFFF;
rommem[17339] <= 16'hFFFF;
rommem[17340] <= 16'hFFFF;
rommem[17341] <= 16'hFFFF;
rommem[17342] <= 16'hFFFF;
rommem[17343] <= 16'hFFFF;
rommem[17344] <= 16'hFFFF;
rommem[17345] <= 16'hFFFF;
rommem[17346] <= 16'hFFFF;
rommem[17347] <= 16'hFFFF;
rommem[17348] <= 16'hFFFF;
rommem[17349] <= 16'hFFFF;
rommem[17350] <= 16'hFFFF;
rommem[17351] <= 16'hFFFF;
rommem[17352] <= 16'hFFFF;
rommem[17353] <= 16'hFFFF;
rommem[17354] <= 16'hFFFF;
rommem[17355] <= 16'hFFFF;
rommem[17356] <= 16'hFFFF;
rommem[17357] <= 16'hFFFF;
rommem[17358] <= 16'hFFFF;
rommem[17359] <= 16'hFFFF;
rommem[17360] <= 16'hFFFF;
rommem[17361] <= 16'hFFFF;
rommem[17362] <= 16'hFFFF;
rommem[17363] <= 16'hFFFF;
rommem[17364] <= 16'hFFFF;
rommem[17365] <= 16'hFFFF;
rommem[17366] <= 16'hFFFF;
rommem[17367] <= 16'hFFFF;
rommem[17368] <= 16'hFFFF;
rommem[17369] <= 16'hFFFF;
rommem[17370] <= 16'hFFFF;
rommem[17371] <= 16'hFFFF;
rommem[17372] <= 16'hFFFF;
rommem[17373] <= 16'hFFFF;
rommem[17374] <= 16'hFFFF;
rommem[17375] <= 16'hFFFF;
rommem[17376] <= 16'hFFFF;
rommem[17377] <= 16'hFFFF;
rommem[17378] <= 16'hFFFF;
rommem[17379] <= 16'hFFFF;
rommem[17380] <= 16'hFFFF;
rommem[17381] <= 16'hFFFF;
rommem[17382] <= 16'hFFFF;
rommem[17383] <= 16'hFFFF;
rommem[17384] <= 16'hFFFF;
rommem[17385] <= 16'hFFFF;
rommem[17386] <= 16'hFFFF;
rommem[17387] <= 16'hFFFF;
rommem[17388] <= 16'hFFFF;
rommem[17389] <= 16'hFFFF;
rommem[17390] <= 16'hFFFF;
rommem[17391] <= 16'hFFFF;
rommem[17392] <= 16'hFFFF;
rommem[17393] <= 16'hFFFF;
rommem[17394] <= 16'hFFFF;
rommem[17395] <= 16'hFFFF;
rommem[17396] <= 16'hFFFF;
rommem[17397] <= 16'hFFFF;
rommem[17398] <= 16'hFFFF;
rommem[17399] <= 16'hFFFF;
rommem[17400] <= 16'hFFFF;
rommem[17401] <= 16'hFFFF;
rommem[17402] <= 16'hFFFF;
rommem[17403] <= 16'hFFFF;
rommem[17404] <= 16'hFFFF;
rommem[17405] <= 16'hFFFF;
rommem[17406] <= 16'hFFFF;
rommem[17407] <= 16'hFFFF;
rommem[17408] <= 16'hFFFF;
rommem[17409] <= 16'hFFFF;
rommem[17410] <= 16'hFFFF;
rommem[17411] <= 16'hFFFF;
rommem[17412] <= 16'hFFFF;
rommem[17413] <= 16'hFFFF;
rommem[17414] <= 16'hFFFF;
rommem[17415] <= 16'hFFFF;
rommem[17416] <= 16'hFFFF;
rommem[17417] <= 16'hFFFF;
rommem[17418] <= 16'hFFFF;
rommem[17419] <= 16'hFFFF;
rommem[17420] <= 16'hFFFF;
rommem[17421] <= 16'hFFFF;
rommem[17422] <= 16'hFFFF;
rommem[17423] <= 16'hFFFF;
rommem[17424] <= 16'hFFFF;
rommem[17425] <= 16'hFFFF;
rommem[17426] <= 16'hFFFF;
rommem[17427] <= 16'hFFFF;
rommem[17428] <= 16'hFFFF;
rommem[17429] <= 16'hFFFF;
rommem[17430] <= 16'hFFFF;
rommem[17431] <= 16'hFFFF;
rommem[17432] <= 16'hFFFF;
rommem[17433] <= 16'hFFFF;
rommem[17434] <= 16'hFFFF;
rommem[17435] <= 16'hFFFF;
rommem[17436] <= 16'hFFFF;
rommem[17437] <= 16'hFFFF;
rommem[17438] <= 16'hFFFF;
rommem[17439] <= 16'hFFFF;
rommem[17440] <= 16'hFFFF;
rommem[17441] <= 16'hFFFF;
rommem[17442] <= 16'hFFFF;
rommem[17443] <= 16'hFFFF;
rommem[17444] <= 16'hFFFF;
rommem[17445] <= 16'hFFFF;
rommem[17446] <= 16'hFFFF;
rommem[17447] <= 16'hFFFF;
rommem[17448] <= 16'hFFFF;
rommem[17449] <= 16'hFFFF;
rommem[17450] <= 16'hFFFF;
rommem[17451] <= 16'hFFFF;
rommem[17452] <= 16'hFFFF;
rommem[17453] <= 16'hFFFF;
rommem[17454] <= 16'hFFFF;
rommem[17455] <= 16'hFFFF;
rommem[17456] <= 16'hFFFF;
rommem[17457] <= 16'hFFFF;
rommem[17458] <= 16'hFFFF;
rommem[17459] <= 16'hFFFF;
rommem[17460] <= 16'hFFFF;
rommem[17461] <= 16'hFFFF;
rommem[17462] <= 16'hFFFF;
rommem[17463] <= 16'hFFFF;
rommem[17464] <= 16'hFFFF;
rommem[17465] <= 16'hFFFF;
rommem[17466] <= 16'hFFFF;
rommem[17467] <= 16'hFFFF;
rommem[17468] <= 16'hFFFF;
rommem[17469] <= 16'hFFFF;
rommem[17470] <= 16'hFFFF;
rommem[17471] <= 16'hFFFF;
rommem[17472] <= 16'hFFFF;
rommem[17473] <= 16'hFFFF;
rommem[17474] <= 16'hFFFF;
rommem[17475] <= 16'hFFFF;
rommem[17476] <= 16'hFFFF;
rommem[17477] <= 16'hFFFF;
rommem[17478] <= 16'hFFFF;
rommem[17479] <= 16'hFFFF;
rommem[17480] <= 16'hFFFF;
rommem[17481] <= 16'hFFFF;
rommem[17482] <= 16'hFFFF;
rommem[17483] <= 16'hFFFF;
rommem[17484] <= 16'hFFFF;
rommem[17485] <= 16'hFFFF;
rommem[17486] <= 16'hFFFF;
rommem[17487] <= 16'hFFFF;
rommem[17488] <= 16'hFFFF;
rommem[17489] <= 16'hFFFF;
rommem[17490] <= 16'hFFFF;
rommem[17491] <= 16'hFFFF;
rommem[17492] <= 16'hFFFF;
rommem[17493] <= 16'hFFFF;
rommem[17494] <= 16'hFFFF;
rommem[17495] <= 16'hFFFF;
rommem[17496] <= 16'hFFFF;
rommem[17497] <= 16'hFFFF;
rommem[17498] <= 16'hFFFF;
rommem[17499] <= 16'hFFFF;
rommem[17500] <= 16'hFFFF;
rommem[17501] <= 16'hFFFF;
rommem[17502] <= 16'hFFFF;
rommem[17503] <= 16'hFFFF;
rommem[17504] <= 16'hFFFF;
rommem[17505] <= 16'hFFFF;
rommem[17506] <= 16'hFFFF;
rommem[17507] <= 16'hFFFF;
rommem[17508] <= 16'hFFFF;
rommem[17509] <= 16'hFFFF;
rommem[17510] <= 16'hFFFF;
rommem[17511] <= 16'hFFFF;
rommem[17512] <= 16'hFFFF;
rommem[17513] <= 16'hFFFF;
rommem[17514] <= 16'hFFFF;
rommem[17515] <= 16'hFFFF;
rommem[17516] <= 16'hFFFF;
rommem[17517] <= 16'hFFFF;
rommem[17518] <= 16'hFFFF;
rommem[17519] <= 16'hFFFF;
rommem[17520] <= 16'hFFFF;
rommem[17521] <= 16'hFFFF;
rommem[17522] <= 16'hFFFF;
rommem[17523] <= 16'hFFFF;
rommem[17524] <= 16'hFFFF;
rommem[17525] <= 16'hFFFF;
rommem[17526] <= 16'hFFFF;
rommem[17527] <= 16'hFFFF;
rommem[17528] <= 16'hFFFF;
rommem[17529] <= 16'hFFFF;
rommem[17530] <= 16'hFFFF;
rommem[17531] <= 16'hFFFF;
rommem[17532] <= 16'hFFFF;
rommem[17533] <= 16'hFFFF;
rommem[17534] <= 16'hFFFF;
rommem[17535] <= 16'hFFFF;
rommem[17536] <= 16'hFFFF;
rommem[17537] <= 16'hFFFF;
rommem[17538] <= 16'hFFFF;
rommem[17539] <= 16'hFFFF;
rommem[17540] <= 16'hFFFF;
rommem[17541] <= 16'hFFFF;
rommem[17542] <= 16'hFFFF;
rommem[17543] <= 16'hFFFF;
rommem[17544] <= 16'hFFFF;
rommem[17545] <= 16'hFFFF;
rommem[17546] <= 16'hFFFF;
rommem[17547] <= 16'hFFFF;
rommem[17548] <= 16'hFFFF;
rommem[17549] <= 16'hFFFF;
rommem[17550] <= 16'hFFFF;
rommem[17551] <= 16'hFFFF;
rommem[17552] <= 16'hFFFF;
rommem[17553] <= 16'hFFFF;
rommem[17554] <= 16'hFFFF;
rommem[17555] <= 16'hFFFF;
rommem[17556] <= 16'hFFFF;
rommem[17557] <= 16'hFFFF;
rommem[17558] <= 16'hFFFF;
rommem[17559] <= 16'hFFFF;
rommem[17560] <= 16'hFFFF;
rommem[17561] <= 16'hFFFF;
rommem[17562] <= 16'hFFFF;
rommem[17563] <= 16'hFFFF;
rommem[17564] <= 16'hFFFF;
rommem[17565] <= 16'hFFFF;
rommem[17566] <= 16'hFFFF;
rommem[17567] <= 16'hFFFF;
rommem[17568] <= 16'hFFFF;
rommem[17569] <= 16'hFFFF;
rommem[17570] <= 16'hFFFF;
rommem[17571] <= 16'hFFFF;
rommem[17572] <= 16'hFFFF;
rommem[17573] <= 16'hFFFF;
rommem[17574] <= 16'hFFFF;
rommem[17575] <= 16'hFFFF;
rommem[17576] <= 16'hFFFF;
rommem[17577] <= 16'hFFFF;
rommem[17578] <= 16'hFFFF;
rommem[17579] <= 16'hFFFF;
rommem[17580] <= 16'hFFFF;
rommem[17581] <= 16'hFFFF;
rommem[17582] <= 16'hFFFF;
rommem[17583] <= 16'hFFFF;
rommem[17584] <= 16'hFFFF;
rommem[17585] <= 16'hFFFF;
rommem[17586] <= 16'hFFFF;
rommem[17587] <= 16'hFFFF;
rommem[17588] <= 16'hFFFF;
rommem[17589] <= 16'hFFFF;
rommem[17590] <= 16'hFFFF;
rommem[17591] <= 16'hFFFF;
rommem[17592] <= 16'hFFFF;
rommem[17593] <= 16'hFFFF;
rommem[17594] <= 16'hFFFF;
rommem[17595] <= 16'hFFFF;
rommem[17596] <= 16'hFFFF;
rommem[17597] <= 16'hFFFF;
rommem[17598] <= 16'hFFFF;
rommem[17599] <= 16'hFFFF;
rommem[17600] <= 16'hFFFF;
rommem[17601] <= 16'hFFFF;
rommem[17602] <= 16'hFFFF;
rommem[17603] <= 16'hFFFF;
rommem[17604] <= 16'hFFFF;
rommem[17605] <= 16'hFFFF;
rommem[17606] <= 16'hFFFF;
rommem[17607] <= 16'hFFFF;
rommem[17608] <= 16'hFFFF;
rommem[17609] <= 16'hFFFF;
rommem[17610] <= 16'hFFFF;
rommem[17611] <= 16'hFFFF;
rommem[17612] <= 16'hFFFF;
rommem[17613] <= 16'hFFFF;
rommem[17614] <= 16'hFFFF;
rommem[17615] <= 16'hFFFF;
rommem[17616] <= 16'hFFFF;
rommem[17617] <= 16'hFFFF;
rommem[17618] <= 16'hFFFF;
rommem[17619] <= 16'hFFFF;
rommem[17620] <= 16'hFFFF;
rommem[17621] <= 16'hFFFF;
rommem[17622] <= 16'hFFFF;
rommem[17623] <= 16'hFFFF;
rommem[17624] <= 16'hFFFF;
rommem[17625] <= 16'hFFFF;
rommem[17626] <= 16'hFFFF;
rommem[17627] <= 16'hFFFF;
rommem[17628] <= 16'hFFFF;
rommem[17629] <= 16'hFFFF;
rommem[17630] <= 16'hFFFF;
rommem[17631] <= 16'hFFFF;
rommem[17632] <= 16'hFFFF;
rommem[17633] <= 16'hFFFF;
rommem[17634] <= 16'hFFFF;
rommem[17635] <= 16'hFFFF;
rommem[17636] <= 16'hFFFF;
rommem[17637] <= 16'hFFFF;
rommem[17638] <= 16'hFFFF;
rommem[17639] <= 16'hFFFF;
rommem[17640] <= 16'hFFFF;
rommem[17641] <= 16'hFFFF;
rommem[17642] <= 16'hFFFF;
rommem[17643] <= 16'hFFFF;
rommem[17644] <= 16'hFFFF;
rommem[17645] <= 16'hFFFF;
rommem[17646] <= 16'hFFFF;
rommem[17647] <= 16'hFFFF;
rommem[17648] <= 16'hFFFF;
rommem[17649] <= 16'hFFFF;
rommem[17650] <= 16'hFFFF;
rommem[17651] <= 16'hFFFF;
rommem[17652] <= 16'hFFFF;
rommem[17653] <= 16'hFFFF;
rommem[17654] <= 16'hFFFF;
rommem[17655] <= 16'hFFFF;
rommem[17656] <= 16'hFFFF;
rommem[17657] <= 16'hFFFF;
rommem[17658] <= 16'hFFFF;
rommem[17659] <= 16'hFFFF;
rommem[17660] <= 16'hFFFF;
rommem[17661] <= 16'hFFFF;
rommem[17662] <= 16'hFFFF;
rommem[17663] <= 16'hFFFF;
rommem[17664] <= 16'hFFFF;
rommem[17665] <= 16'hFFFF;
rommem[17666] <= 16'hFFFF;
rommem[17667] <= 16'hFFFF;
rommem[17668] <= 16'hFFFF;
rommem[17669] <= 16'hFFFF;
rommem[17670] <= 16'hFFFF;
rommem[17671] <= 16'hFFFF;
rommem[17672] <= 16'hFFFF;
rommem[17673] <= 16'hFFFF;
rommem[17674] <= 16'hFFFF;
rommem[17675] <= 16'hFFFF;
rommem[17676] <= 16'hFFFF;
rommem[17677] <= 16'hFFFF;
rommem[17678] <= 16'hFFFF;
rommem[17679] <= 16'hFFFF;
rommem[17680] <= 16'hFFFF;
rommem[17681] <= 16'hFFFF;
rommem[17682] <= 16'hFFFF;
rommem[17683] <= 16'hFFFF;
rommem[17684] <= 16'hFFFF;
rommem[17685] <= 16'hFFFF;
rommem[17686] <= 16'hFFFF;
rommem[17687] <= 16'hFFFF;
rommem[17688] <= 16'hFFFF;
rommem[17689] <= 16'hFFFF;
rommem[17690] <= 16'hFFFF;
rommem[17691] <= 16'hFFFF;
rommem[17692] <= 16'hFFFF;
rommem[17693] <= 16'hFFFF;
rommem[17694] <= 16'hFFFF;
rommem[17695] <= 16'hFFFF;
rommem[17696] <= 16'hFFFF;
rommem[17697] <= 16'hFFFF;
rommem[17698] <= 16'hFFFF;
rommem[17699] <= 16'hFFFF;
rommem[17700] <= 16'hFFFF;
rommem[17701] <= 16'hFFFF;
rommem[17702] <= 16'hFFFF;
rommem[17703] <= 16'hFFFF;
rommem[17704] <= 16'hFFFF;
rommem[17705] <= 16'hFFFF;
rommem[17706] <= 16'hFFFF;
rommem[17707] <= 16'hFFFF;
rommem[17708] <= 16'hFFFF;
rommem[17709] <= 16'hFFFF;
rommem[17710] <= 16'hFFFF;
rommem[17711] <= 16'hFFFF;
rommem[17712] <= 16'hFFFF;
rommem[17713] <= 16'hFFFF;
rommem[17714] <= 16'hFFFF;
rommem[17715] <= 16'hFFFF;
rommem[17716] <= 16'hFFFF;
rommem[17717] <= 16'hFFFF;
rommem[17718] <= 16'hFFFF;
rommem[17719] <= 16'hFFFF;
rommem[17720] <= 16'hFFFF;
rommem[17721] <= 16'hFFFF;
rommem[17722] <= 16'hFFFF;
rommem[17723] <= 16'hFFFF;
rommem[17724] <= 16'hFFFF;
rommem[17725] <= 16'hFFFF;
rommem[17726] <= 16'hFFFF;
rommem[17727] <= 16'hFFFF;
rommem[17728] <= 16'hFFFF;
rommem[17729] <= 16'hFFFF;
rommem[17730] <= 16'hFFFF;
rommem[17731] <= 16'hFFFF;
rommem[17732] <= 16'hFFFF;
rommem[17733] <= 16'hFFFF;
rommem[17734] <= 16'hFFFF;
rommem[17735] <= 16'hFFFF;
rommem[17736] <= 16'hFFFF;
rommem[17737] <= 16'hFFFF;
rommem[17738] <= 16'hFFFF;
rommem[17739] <= 16'hFFFF;
rommem[17740] <= 16'hFFFF;
rommem[17741] <= 16'hFFFF;
rommem[17742] <= 16'hFFFF;
rommem[17743] <= 16'hFFFF;
rommem[17744] <= 16'hFFFF;
rommem[17745] <= 16'hFFFF;
rommem[17746] <= 16'hFFFF;
rommem[17747] <= 16'hFFFF;
rommem[17748] <= 16'hFFFF;
rommem[17749] <= 16'hFFFF;
rommem[17750] <= 16'hFFFF;
rommem[17751] <= 16'hFFFF;
rommem[17752] <= 16'hFFFF;
rommem[17753] <= 16'hFFFF;
rommem[17754] <= 16'hFFFF;
rommem[17755] <= 16'hFFFF;
rommem[17756] <= 16'hFFFF;
rommem[17757] <= 16'hFFFF;
rommem[17758] <= 16'hFFFF;
rommem[17759] <= 16'hFFFF;
rommem[17760] <= 16'hFFFF;
rommem[17761] <= 16'hFFFF;
rommem[17762] <= 16'hFFFF;
rommem[17763] <= 16'hFFFF;
rommem[17764] <= 16'hFFFF;
rommem[17765] <= 16'hFFFF;
rommem[17766] <= 16'hFFFF;
rommem[17767] <= 16'hFFFF;
rommem[17768] <= 16'hFFFF;
rommem[17769] <= 16'hFFFF;
rommem[17770] <= 16'hFFFF;
rommem[17771] <= 16'hFFFF;
rommem[17772] <= 16'hFFFF;
rommem[17773] <= 16'hFFFF;
rommem[17774] <= 16'hFFFF;
rommem[17775] <= 16'hFFFF;
rommem[17776] <= 16'hFFFF;
rommem[17777] <= 16'hFFFF;
rommem[17778] <= 16'hFFFF;
rommem[17779] <= 16'hFFFF;
rommem[17780] <= 16'hFFFF;
rommem[17781] <= 16'hFFFF;
rommem[17782] <= 16'hFFFF;
rommem[17783] <= 16'hFFFF;
rommem[17784] <= 16'hFFFF;
rommem[17785] <= 16'hFFFF;
rommem[17786] <= 16'hFFFF;
rommem[17787] <= 16'hFFFF;
rommem[17788] <= 16'hFFFF;
rommem[17789] <= 16'hFFFF;
rommem[17790] <= 16'hFFFF;
rommem[17791] <= 16'hFFFF;
rommem[17792] <= 16'hFFFF;
rommem[17793] <= 16'hFFFF;
rommem[17794] <= 16'hFFFF;
rommem[17795] <= 16'hFFFF;
rommem[17796] <= 16'hFFFF;
rommem[17797] <= 16'hFFFF;
rommem[17798] <= 16'hFFFF;
rommem[17799] <= 16'hFFFF;
rommem[17800] <= 16'hFFFF;
rommem[17801] <= 16'hFFFF;
rommem[17802] <= 16'hFFFF;
rommem[17803] <= 16'hFFFF;
rommem[17804] <= 16'hFFFF;
rommem[17805] <= 16'hFFFF;
rommem[17806] <= 16'hFFFF;
rommem[17807] <= 16'hFFFF;
rommem[17808] <= 16'hFFFF;
rommem[17809] <= 16'hFFFF;
rommem[17810] <= 16'hFFFF;
rommem[17811] <= 16'hFFFF;
rommem[17812] <= 16'hFFFF;
rommem[17813] <= 16'hFFFF;
rommem[17814] <= 16'hFFFF;
rommem[17815] <= 16'hFFFF;
rommem[17816] <= 16'hFFFF;
rommem[17817] <= 16'hFFFF;
rommem[17818] <= 16'hFFFF;
rommem[17819] <= 16'hFFFF;
rommem[17820] <= 16'hFFFF;
rommem[17821] <= 16'hFFFF;
rommem[17822] <= 16'hFFFF;
rommem[17823] <= 16'hFFFF;
rommem[17824] <= 16'hFFFF;
rommem[17825] <= 16'hFFFF;
rommem[17826] <= 16'hFFFF;
rommem[17827] <= 16'hFFFF;
rommem[17828] <= 16'hFFFF;
rommem[17829] <= 16'hFFFF;
rommem[17830] <= 16'hFFFF;
rommem[17831] <= 16'hFFFF;
rommem[17832] <= 16'hFFFF;
rommem[17833] <= 16'hFFFF;
rommem[17834] <= 16'hFFFF;
rommem[17835] <= 16'hFFFF;
rommem[17836] <= 16'hFFFF;
rommem[17837] <= 16'hFFFF;
rommem[17838] <= 16'hFFFF;
rommem[17839] <= 16'hFFFF;
rommem[17840] <= 16'hFFFF;
rommem[17841] <= 16'hFFFF;
rommem[17842] <= 16'hFFFF;
rommem[17843] <= 16'hFFFF;
rommem[17844] <= 16'hFFFF;
rommem[17845] <= 16'hFFFF;
rommem[17846] <= 16'hFFFF;
rommem[17847] <= 16'hFFFF;
rommem[17848] <= 16'hFFFF;
rommem[17849] <= 16'hFFFF;
rommem[17850] <= 16'hFFFF;
rommem[17851] <= 16'hFFFF;
rommem[17852] <= 16'hFFFF;
rommem[17853] <= 16'hFFFF;
rommem[17854] <= 16'hFFFF;
rommem[17855] <= 16'hFFFF;
rommem[17856] <= 16'hFFFF;
rommem[17857] <= 16'hFFFF;
rommem[17858] <= 16'hFFFF;
rommem[17859] <= 16'hFFFF;
rommem[17860] <= 16'hFFFF;
rommem[17861] <= 16'hFFFF;
rommem[17862] <= 16'hFFFF;
rommem[17863] <= 16'hFFFF;
rommem[17864] <= 16'hFFFF;
rommem[17865] <= 16'hFFFF;
rommem[17866] <= 16'hFFFF;
rommem[17867] <= 16'hFFFF;
rommem[17868] <= 16'hFFFF;
rommem[17869] <= 16'hFFFF;
rommem[17870] <= 16'hFFFF;
rommem[17871] <= 16'hFFFF;
rommem[17872] <= 16'hFFFF;
rommem[17873] <= 16'hFFFF;
rommem[17874] <= 16'hFFFF;
rommem[17875] <= 16'hFFFF;
rommem[17876] <= 16'hFFFF;
rommem[17877] <= 16'hFFFF;
rommem[17878] <= 16'hFFFF;
rommem[17879] <= 16'hFFFF;
rommem[17880] <= 16'hFFFF;
rommem[17881] <= 16'hFFFF;
rommem[17882] <= 16'hFFFF;
rommem[17883] <= 16'hFFFF;
rommem[17884] <= 16'hFFFF;
rommem[17885] <= 16'hFFFF;
rommem[17886] <= 16'hFFFF;
rommem[17887] <= 16'hFFFF;
rommem[17888] <= 16'hFFFF;
rommem[17889] <= 16'hFFFF;
rommem[17890] <= 16'hFFFF;
rommem[17891] <= 16'hFFFF;
rommem[17892] <= 16'hFFFF;
rommem[17893] <= 16'hFFFF;
rommem[17894] <= 16'hFFFF;
rommem[17895] <= 16'hFFFF;
rommem[17896] <= 16'hFFFF;
rommem[17897] <= 16'hFFFF;
rommem[17898] <= 16'hFFFF;
rommem[17899] <= 16'hFFFF;
rommem[17900] <= 16'hFFFF;
rommem[17901] <= 16'hFFFF;
rommem[17902] <= 16'hFFFF;
rommem[17903] <= 16'hFFFF;
rommem[17904] <= 16'hFFFF;
rommem[17905] <= 16'hFFFF;
rommem[17906] <= 16'hFFFF;
rommem[17907] <= 16'hFFFF;
rommem[17908] <= 16'hFFFF;
rommem[17909] <= 16'hFFFF;
rommem[17910] <= 16'hFFFF;
rommem[17911] <= 16'hFFFF;
rommem[17912] <= 16'hFFFF;
rommem[17913] <= 16'hFFFF;
rommem[17914] <= 16'hFFFF;
rommem[17915] <= 16'hFFFF;
rommem[17916] <= 16'hFFFF;
rommem[17917] <= 16'hFFFF;
rommem[17918] <= 16'hFFFF;
rommem[17919] <= 16'hFFFF;
rommem[17920] <= 16'hFFFF;
rommem[17921] <= 16'hFFFF;
rommem[17922] <= 16'hFFFF;
rommem[17923] <= 16'hFFFF;
rommem[17924] <= 16'hFFFF;
rommem[17925] <= 16'hFFFF;
rommem[17926] <= 16'hFFFF;
rommem[17927] <= 16'hFFFF;
rommem[17928] <= 16'hFFFF;
rommem[17929] <= 16'hFFFF;
rommem[17930] <= 16'hFFFF;
rommem[17931] <= 16'hFFFF;
rommem[17932] <= 16'hFFFF;
rommem[17933] <= 16'hFFFF;
rommem[17934] <= 16'hFFFF;
rommem[17935] <= 16'hFFFF;
rommem[17936] <= 16'hFFFF;
rommem[17937] <= 16'hFFFF;
rommem[17938] <= 16'hFFFF;
rommem[17939] <= 16'hFFFF;
rommem[17940] <= 16'hFFFF;
rommem[17941] <= 16'hFFFF;
rommem[17942] <= 16'hFFFF;
rommem[17943] <= 16'hFFFF;
rommem[17944] <= 16'hFFFF;
rommem[17945] <= 16'hFFFF;
rommem[17946] <= 16'hFFFF;
rommem[17947] <= 16'hFFFF;
rommem[17948] <= 16'hFFFF;
rommem[17949] <= 16'hFFFF;
rommem[17950] <= 16'hFFFF;
rommem[17951] <= 16'hFFFF;
rommem[17952] <= 16'hFFFF;
rommem[17953] <= 16'hFFFF;
rommem[17954] <= 16'hFFFF;
rommem[17955] <= 16'hFFFF;
rommem[17956] <= 16'hFFFF;
rommem[17957] <= 16'hFFFF;
rommem[17958] <= 16'hFFFF;
rommem[17959] <= 16'hFFFF;
rommem[17960] <= 16'hFFFF;
rommem[17961] <= 16'hFFFF;
rommem[17962] <= 16'hFFFF;
rommem[17963] <= 16'hFFFF;
rommem[17964] <= 16'hFFFF;
rommem[17965] <= 16'hFFFF;
rommem[17966] <= 16'hFFFF;
rommem[17967] <= 16'hFFFF;
rommem[17968] <= 16'hFFFF;
rommem[17969] <= 16'hFFFF;
rommem[17970] <= 16'hFFFF;
rommem[17971] <= 16'hFFFF;
rommem[17972] <= 16'hFFFF;
rommem[17973] <= 16'hFFFF;
rommem[17974] <= 16'hFFFF;
rommem[17975] <= 16'hFFFF;
rommem[17976] <= 16'hFFFF;
rommem[17977] <= 16'hFFFF;
rommem[17978] <= 16'hFFFF;
rommem[17979] <= 16'hFFFF;
rommem[17980] <= 16'hFFFF;
rommem[17981] <= 16'hFFFF;
rommem[17982] <= 16'hFFFF;
rommem[17983] <= 16'hFFFF;
rommem[17984] <= 16'hFFFF;
rommem[17985] <= 16'hFFFF;
rommem[17986] <= 16'hFFFF;
rommem[17987] <= 16'hFFFF;
rommem[17988] <= 16'hFFFF;
rommem[17989] <= 16'hFFFF;
rommem[17990] <= 16'hFFFF;
rommem[17991] <= 16'hFFFF;
rommem[17992] <= 16'hFFFF;
rommem[17993] <= 16'hFFFF;
rommem[17994] <= 16'hFFFF;
rommem[17995] <= 16'hFFFF;
rommem[17996] <= 16'hFFFF;
rommem[17997] <= 16'hFFFF;
rommem[17998] <= 16'hFFFF;
rommem[17999] <= 16'hFFFF;
rommem[18000] <= 16'hFFFF;
rommem[18001] <= 16'hFFFF;
rommem[18002] <= 16'hFFFF;
rommem[18003] <= 16'hFFFF;
rommem[18004] <= 16'hFFFF;
rommem[18005] <= 16'hFFFF;
rommem[18006] <= 16'hFFFF;
rommem[18007] <= 16'hFFFF;
rommem[18008] <= 16'hFFFF;
rommem[18009] <= 16'hFFFF;
rommem[18010] <= 16'hFFFF;
rommem[18011] <= 16'hFFFF;
rommem[18012] <= 16'hFFFF;
rommem[18013] <= 16'hFFFF;
rommem[18014] <= 16'hFFFF;
rommem[18015] <= 16'hFFFF;
rommem[18016] <= 16'hFFFF;
rommem[18017] <= 16'hFFFF;
rommem[18018] <= 16'hFFFF;
rommem[18019] <= 16'hFFFF;
rommem[18020] <= 16'hFFFF;
rommem[18021] <= 16'hFFFF;
rommem[18022] <= 16'hFFFF;
rommem[18023] <= 16'hFFFF;
rommem[18024] <= 16'hFFFF;
rommem[18025] <= 16'hFFFF;
rommem[18026] <= 16'hFFFF;
rommem[18027] <= 16'hFFFF;
rommem[18028] <= 16'hFFFF;
rommem[18029] <= 16'hFFFF;
rommem[18030] <= 16'hFFFF;
rommem[18031] <= 16'hFFFF;
rommem[18032] <= 16'hFFFF;
rommem[18033] <= 16'hFFFF;
rommem[18034] <= 16'hFFFF;
rommem[18035] <= 16'hFFFF;
rommem[18036] <= 16'hFFFF;
rommem[18037] <= 16'hFFFF;
rommem[18038] <= 16'hFFFF;
rommem[18039] <= 16'hFFFF;
rommem[18040] <= 16'hFFFF;
rommem[18041] <= 16'hFFFF;
rommem[18042] <= 16'hFFFF;
rommem[18043] <= 16'hFFFF;
rommem[18044] <= 16'hFFFF;
rommem[18045] <= 16'hFFFF;
rommem[18046] <= 16'hFFFF;
rommem[18047] <= 16'hFFFF;
rommem[18048] <= 16'hFFFF;
rommem[18049] <= 16'hFFFF;
rommem[18050] <= 16'hFFFF;
rommem[18051] <= 16'hFFFF;
rommem[18052] <= 16'hFFFF;
rommem[18053] <= 16'hFFFF;
rommem[18054] <= 16'hFFFF;
rommem[18055] <= 16'hFFFF;
rommem[18056] <= 16'hFFFF;
rommem[18057] <= 16'hFFFF;
rommem[18058] <= 16'hFFFF;
rommem[18059] <= 16'hFFFF;
rommem[18060] <= 16'hFFFF;
rommem[18061] <= 16'hFFFF;
rommem[18062] <= 16'hFFFF;
rommem[18063] <= 16'hFFFF;
rommem[18064] <= 16'hFFFF;
rommem[18065] <= 16'hFFFF;
rommem[18066] <= 16'hFFFF;
rommem[18067] <= 16'hFFFF;
rommem[18068] <= 16'hFFFF;
rommem[18069] <= 16'hFFFF;
rommem[18070] <= 16'hFFFF;
rommem[18071] <= 16'hFFFF;
rommem[18072] <= 16'hFFFF;
rommem[18073] <= 16'hFFFF;
rommem[18074] <= 16'hFFFF;
rommem[18075] <= 16'hFFFF;
rommem[18076] <= 16'hFFFF;
rommem[18077] <= 16'hFFFF;
rommem[18078] <= 16'hFFFF;
rommem[18079] <= 16'hFFFF;
rommem[18080] <= 16'hFFFF;
rommem[18081] <= 16'hFFFF;
rommem[18082] <= 16'hFFFF;
rommem[18083] <= 16'hFFFF;
rommem[18084] <= 16'hFFFF;
rommem[18085] <= 16'hFFFF;
rommem[18086] <= 16'hFFFF;
rommem[18087] <= 16'hFFFF;
rommem[18088] <= 16'hFFFF;
rommem[18089] <= 16'hFFFF;
rommem[18090] <= 16'hFFFF;
rommem[18091] <= 16'hFFFF;
rommem[18092] <= 16'hFFFF;
rommem[18093] <= 16'hFFFF;
rommem[18094] <= 16'hFFFF;
rommem[18095] <= 16'hFFFF;
rommem[18096] <= 16'hFFFF;
rommem[18097] <= 16'hFFFF;
rommem[18098] <= 16'hFFFF;
rommem[18099] <= 16'hFFFF;
rommem[18100] <= 16'hFFFF;
rommem[18101] <= 16'hFFFF;
rommem[18102] <= 16'hFFFF;
rommem[18103] <= 16'hFFFF;
rommem[18104] <= 16'hFFFF;
rommem[18105] <= 16'hFFFF;
rommem[18106] <= 16'hFFFF;
rommem[18107] <= 16'hFFFF;
rommem[18108] <= 16'hFFFF;
rommem[18109] <= 16'hFFFF;
rommem[18110] <= 16'hFFFF;
rommem[18111] <= 16'hFFFF;
rommem[18112] <= 16'hFFFF;
rommem[18113] <= 16'hFFFF;
rommem[18114] <= 16'hFFFF;
rommem[18115] <= 16'hFFFF;
rommem[18116] <= 16'hFFFF;
rommem[18117] <= 16'hFFFF;
rommem[18118] <= 16'hFFFF;
rommem[18119] <= 16'hFFFF;
rommem[18120] <= 16'hFFFF;
rommem[18121] <= 16'hFFFF;
rommem[18122] <= 16'hFFFF;
rommem[18123] <= 16'hFFFF;
rommem[18124] <= 16'hFFFF;
rommem[18125] <= 16'hFFFF;
rommem[18126] <= 16'hFFFF;
rommem[18127] <= 16'hFFFF;
rommem[18128] <= 16'hFFFF;
rommem[18129] <= 16'hFFFF;
rommem[18130] <= 16'hFFFF;
rommem[18131] <= 16'hFFFF;
rommem[18132] <= 16'hFFFF;
rommem[18133] <= 16'hFFFF;
rommem[18134] <= 16'hFFFF;
rommem[18135] <= 16'hFFFF;
rommem[18136] <= 16'hFFFF;
rommem[18137] <= 16'hFFFF;
rommem[18138] <= 16'hFFFF;
rommem[18139] <= 16'hFFFF;
rommem[18140] <= 16'hFFFF;
rommem[18141] <= 16'hFFFF;
rommem[18142] <= 16'hFFFF;
rommem[18143] <= 16'hFFFF;
rommem[18144] <= 16'hFFFF;
rommem[18145] <= 16'hFFFF;
rommem[18146] <= 16'hFFFF;
rommem[18147] <= 16'hFFFF;
rommem[18148] <= 16'hFFFF;
rommem[18149] <= 16'hFFFF;
rommem[18150] <= 16'hFFFF;
rommem[18151] <= 16'hFFFF;
rommem[18152] <= 16'hFFFF;
rommem[18153] <= 16'hFFFF;
rommem[18154] <= 16'hFFFF;
rommem[18155] <= 16'hFFFF;
rommem[18156] <= 16'hFFFF;
rommem[18157] <= 16'hFFFF;
rommem[18158] <= 16'hFFFF;
rommem[18159] <= 16'hFFFF;
rommem[18160] <= 16'hFFFF;
rommem[18161] <= 16'hFFFF;
rommem[18162] <= 16'hFFFF;
rommem[18163] <= 16'hFFFF;
rommem[18164] <= 16'hFFFF;
rommem[18165] <= 16'hFFFF;
rommem[18166] <= 16'hFFFF;
rommem[18167] <= 16'hFFFF;
rommem[18168] <= 16'hFFFF;
rommem[18169] <= 16'hFFFF;
rommem[18170] <= 16'hFFFF;
rommem[18171] <= 16'hFFFF;
rommem[18172] <= 16'hFFFF;
rommem[18173] <= 16'hFFFF;
rommem[18174] <= 16'hFFFF;
rommem[18175] <= 16'hFFFF;
rommem[18176] <= 16'hFFFF;
rommem[18177] <= 16'hFFFF;
rommem[18178] <= 16'hFFFF;
rommem[18179] <= 16'hFFFF;
rommem[18180] <= 16'hFFFF;
rommem[18181] <= 16'hFFFF;
rommem[18182] <= 16'hFFFF;
rommem[18183] <= 16'hFFFF;
rommem[18184] <= 16'hFFFF;
rommem[18185] <= 16'hFFFF;
rommem[18186] <= 16'hFFFF;
rommem[18187] <= 16'hFFFF;
rommem[18188] <= 16'hFFFF;
rommem[18189] <= 16'hFFFF;
rommem[18190] <= 16'hFFFF;
rommem[18191] <= 16'hFFFF;
rommem[18192] <= 16'hFFFF;
rommem[18193] <= 16'hFFFF;
rommem[18194] <= 16'hFFFF;
rommem[18195] <= 16'hFFFF;
rommem[18196] <= 16'hFFFF;
rommem[18197] <= 16'hFFFF;
rommem[18198] <= 16'hFFFF;
rommem[18199] <= 16'hFFFF;
rommem[18200] <= 16'hFFFF;
rommem[18201] <= 16'hFFFF;
rommem[18202] <= 16'hFFFF;
rommem[18203] <= 16'hFFFF;
rommem[18204] <= 16'hFFFF;
rommem[18205] <= 16'hFFFF;
rommem[18206] <= 16'hFFFF;
rommem[18207] <= 16'hFFFF;
rommem[18208] <= 16'hFFFF;
rommem[18209] <= 16'hFFFF;
rommem[18210] <= 16'hFFFF;
rommem[18211] <= 16'hFFFF;
rommem[18212] <= 16'hFFFF;
rommem[18213] <= 16'hFFFF;
rommem[18214] <= 16'hFFFF;
rommem[18215] <= 16'hFFFF;
rommem[18216] <= 16'hFFFF;
rommem[18217] <= 16'hFFFF;
rommem[18218] <= 16'hFFFF;
rommem[18219] <= 16'hFFFF;
rommem[18220] <= 16'hFFFF;
rommem[18221] <= 16'hFFFF;
rommem[18222] <= 16'hFFFF;
rommem[18223] <= 16'hFFFF;
rommem[18224] <= 16'hFFFF;
rommem[18225] <= 16'hFFFF;
rommem[18226] <= 16'hFFFF;
rommem[18227] <= 16'hFFFF;
rommem[18228] <= 16'hFFFF;
rommem[18229] <= 16'hFFFF;
rommem[18230] <= 16'hFFFF;
rommem[18231] <= 16'hFFFF;
rommem[18232] <= 16'hFFFF;
rommem[18233] <= 16'hFFFF;
rommem[18234] <= 16'hFFFF;
rommem[18235] <= 16'hFFFF;
rommem[18236] <= 16'hFFFF;
rommem[18237] <= 16'hFFFF;
rommem[18238] <= 16'hFFFF;
rommem[18239] <= 16'hFFFF;
rommem[18240] <= 16'hFFFF;
rommem[18241] <= 16'hFFFF;
rommem[18242] <= 16'hFFFF;
rommem[18243] <= 16'hFFFF;
rommem[18244] <= 16'hFFFF;
rommem[18245] <= 16'hFFFF;
rommem[18246] <= 16'hFFFF;
rommem[18247] <= 16'hFFFF;
rommem[18248] <= 16'hFFFF;
rommem[18249] <= 16'hFFFF;
rommem[18250] <= 16'hFFFF;
rommem[18251] <= 16'hFFFF;
rommem[18252] <= 16'hFFFF;
rommem[18253] <= 16'hFFFF;
rommem[18254] <= 16'hFFFF;
rommem[18255] <= 16'hFFFF;
rommem[18256] <= 16'hFFFF;
rommem[18257] <= 16'hFFFF;
rommem[18258] <= 16'hFFFF;
rommem[18259] <= 16'hFFFF;
rommem[18260] <= 16'hFFFF;
rommem[18261] <= 16'hFFFF;
rommem[18262] <= 16'hFFFF;
rommem[18263] <= 16'hFFFF;
rommem[18264] <= 16'hFFFF;
rommem[18265] <= 16'hFFFF;
rommem[18266] <= 16'hFFFF;
rommem[18267] <= 16'hFFFF;
rommem[18268] <= 16'hFFFF;
rommem[18269] <= 16'hFFFF;
rommem[18270] <= 16'hFFFF;
rommem[18271] <= 16'hFFFF;
rommem[18272] <= 16'hFFFF;
rommem[18273] <= 16'hFFFF;
rommem[18274] <= 16'hFFFF;
rommem[18275] <= 16'hFFFF;
rommem[18276] <= 16'hFFFF;
rommem[18277] <= 16'hFFFF;
rommem[18278] <= 16'hFFFF;
rommem[18279] <= 16'hFFFF;
rommem[18280] <= 16'hFFFF;
rommem[18281] <= 16'hFFFF;
rommem[18282] <= 16'hFFFF;
rommem[18283] <= 16'hFFFF;
rommem[18284] <= 16'hFFFF;
rommem[18285] <= 16'hFFFF;
rommem[18286] <= 16'hFFFF;
rommem[18287] <= 16'hFFFF;
rommem[18288] <= 16'hFFFF;
rommem[18289] <= 16'hFFFF;
rommem[18290] <= 16'hFFFF;
rommem[18291] <= 16'hFFFF;
rommem[18292] <= 16'hFFFF;
rommem[18293] <= 16'hFFFF;
rommem[18294] <= 16'hFFFF;
rommem[18295] <= 16'hFFFF;
rommem[18296] <= 16'hFFFF;
rommem[18297] <= 16'hFFFF;
rommem[18298] <= 16'hFFFF;
rommem[18299] <= 16'hFFFF;
rommem[18300] <= 16'hFFFF;
rommem[18301] <= 16'hFFFF;
rommem[18302] <= 16'hFFFF;
rommem[18303] <= 16'hFFFF;
rommem[18304] <= 16'hFFFF;
rommem[18305] <= 16'hFFFF;
rommem[18306] <= 16'hFFFF;
rommem[18307] <= 16'hFFFF;
rommem[18308] <= 16'hFFFF;
rommem[18309] <= 16'hFFFF;
rommem[18310] <= 16'hFFFF;
rommem[18311] <= 16'hFFFF;
rommem[18312] <= 16'hFFFF;
rommem[18313] <= 16'hFFFF;
rommem[18314] <= 16'hFFFF;
rommem[18315] <= 16'hFFFF;
rommem[18316] <= 16'hFFFF;
rommem[18317] <= 16'hFFFF;
rommem[18318] <= 16'hFFFF;
rommem[18319] <= 16'hFFFF;
rommem[18320] <= 16'hFFFF;
rommem[18321] <= 16'hFFFF;
rommem[18322] <= 16'hFFFF;
rommem[18323] <= 16'hFFFF;
rommem[18324] <= 16'hFFFF;
rommem[18325] <= 16'hFFFF;
rommem[18326] <= 16'hFFFF;
rommem[18327] <= 16'hFFFF;
rommem[18328] <= 16'hFFFF;
rommem[18329] <= 16'hFFFF;
rommem[18330] <= 16'hFFFF;
rommem[18331] <= 16'hFFFF;
rommem[18332] <= 16'hFFFF;
rommem[18333] <= 16'hFFFF;
rommem[18334] <= 16'hFFFF;
rommem[18335] <= 16'hFFFF;
rommem[18336] <= 16'hFFFF;
rommem[18337] <= 16'hFFFF;
rommem[18338] <= 16'hFFFF;
rommem[18339] <= 16'hFFFF;
rommem[18340] <= 16'hFFFF;
rommem[18341] <= 16'hFFFF;
rommem[18342] <= 16'hFFFF;
rommem[18343] <= 16'hFFFF;
rommem[18344] <= 16'hFFFF;
rommem[18345] <= 16'hFFFF;
rommem[18346] <= 16'hFFFF;
rommem[18347] <= 16'hFFFF;
rommem[18348] <= 16'hFFFF;
rommem[18349] <= 16'hFFFF;
rommem[18350] <= 16'hFFFF;
rommem[18351] <= 16'hFFFF;
rommem[18352] <= 16'hFFFF;
rommem[18353] <= 16'hFFFF;
rommem[18354] <= 16'hFFFF;
rommem[18355] <= 16'hFFFF;
rommem[18356] <= 16'hFFFF;
rommem[18357] <= 16'hFFFF;
rommem[18358] <= 16'hFFFF;
rommem[18359] <= 16'hFFFF;
rommem[18360] <= 16'hFFFF;
rommem[18361] <= 16'hFFFF;
rommem[18362] <= 16'hFFFF;
rommem[18363] <= 16'hFFFF;
rommem[18364] <= 16'hFFFF;
rommem[18365] <= 16'hFFFF;
rommem[18366] <= 16'hFFFF;
rommem[18367] <= 16'hFFFF;
rommem[18368] <= 16'hFFFF;
rommem[18369] <= 16'hFFFF;
rommem[18370] <= 16'hFFFF;
rommem[18371] <= 16'hFFFF;
rommem[18372] <= 16'hFFFF;
rommem[18373] <= 16'hFFFF;
rommem[18374] <= 16'hFFFF;
rommem[18375] <= 16'hFFFF;
rommem[18376] <= 16'hFFFF;
rommem[18377] <= 16'hFFFF;
rommem[18378] <= 16'hFFFF;
rommem[18379] <= 16'hFFFF;
rommem[18380] <= 16'hFFFF;
rommem[18381] <= 16'hFFFF;
rommem[18382] <= 16'hFFFF;
rommem[18383] <= 16'hFFFF;
rommem[18384] <= 16'hFFFF;
rommem[18385] <= 16'hFFFF;
rommem[18386] <= 16'hFFFF;
rommem[18387] <= 16'hFFFF;
rommem[18388] <= 16'hFFFF;
rommem[18389] <= 16'hFFFF;
rommem[18390] <= 16'hFFFF;
rommem[18391] <= 16'hFFFF;
rommem[18392] <= 16'hFFFF;
rommem[18393] <= 16'hFFFF;
rommem[18394] <= 16'hFFFF;
rommem[18395] <= 16'hFFFF;
rommem[18396] <= 16'hFFFF;
rommem[18397] <= 16'hFFFF;
rommem[18398] <= 16'hFFFF;
rommem[18399] <= 16'hFFFF;
rommem[18400] <= 16'hFFFF;
rommem[18401] <= 16'hFFFF;
rommem[18402] <= 16'hFFFF;
rommem[18403] <= 16'hFFFF;
rommem[18404] <= 16'hFFFF;
rommem[18405] <= 16'hFFFF;
rommem[18406] <= 16'hFFFF;
rommem[18407] <= 16'hFFFF;
rommem[18408] <= 16'hFFFF;
rommem[18409] <= 16'hFFFF;
rommem[18410] <= 16'hFFFF;
rommem[18411] <= 16'hFFFF;
rommem[18412] <= 16'hFFFF;
rommem[18413] <= 16'hFFFF;
rommem[18414] <= 16'hFFFF;
rommem[18415] <= 16'hFFFF;
rommem[18416] <= 16'hFFFF;
rommem[18417] <= 16'hFFFF;
rommem[18418] <= 16'hFFFF;
rommem[18419] <= 16'hFFFF;
rommem[18420] <= 16'hFFFF;
rommem[18421] <= 16'hFFFF;
rommem[18422] <= 16'hFFFF;
rommem[18423] <= 16'hFFFF;
rommem[18424] <= 16'hFFFF;
rommem[18425] <= 16'hFFFF;
rommem[18426] <= 16'hFFFF;
rommem[18427] <= 16'hFFFF;
rommem[18428] <= 16'hFFFF;
rommem[18429] <= 16'hFFFF;
rommem[18430] <= 16'hFFFF;
rommem[18431] <= 16'hFFFF;
rommem[18432] <= 16'hFFFF;
rommem[18433] <= 16'hFFFF;
rommem[18434] <= 16'hFFFF;
rommem[18435] <= 16'hFFFF;
rommem[18436] <= 16'hFFFF;
rommem[18437] <= 16'hFFFF;
rommem[18438] <= 16'hFFFF;
rommem[18439] <= 16'hFFFF;
rommem[18440] <= 16'hFFFF;
rommem[18441] <= 16'hFFFF;
rommem[18442] <= 16'hFFFF;
rommem[18443] <= 16'hFFFF;
rommem[18444] <= 16'hFFFF;
rommem[18445] <= 16'hFFFF;
rommem[18446] <= 16'hFFFF;
rommem[18447] <= 16'hFFFF;
rommem[18448] <= 16'hFFFF;
rommem[18449] <= 16'hFFFF;
rommem[18450] <= 16'hFFFF;
rommem[18451] <= 16'hFFFF;
rommem[18452] <= 16'hFFFF;
rommem[18453] <= 16'hFFFF;
rommem[18454] <= 16'hFFFF;
rommem[18455] <= 16'hFFFF;
rommem[18456] <= 16'hFFFF;
rommem[18457] <= 16'hFFFF;
rommem[18458] <= 16'hFFFF;
rommem[18459] <= 16'hFFFF;
rommem[18460] <= 16'hFFFF;
rommem[18461] <= 16'hFFFF;
rommem[18462] <= 16'hFFFF;
rommem[18463] <= 16'hFFFF;
rommem[18464] <= 16'hFFFF;
rommem[18465] <= 16'hFFFF;
rommem[18466] <= 16'hFFFF;
rommem[18467] <= 16'hFFFF;
rommem[18468] <= 16'hFFFF;
rommem[18469] <= 16'hFFFF;
rommem[18470] <= 16'hFFFF;
rommem[18471] <= 16'hFFFF;
rommem[18472] <= 16'hFFFF;
rommem[18473] <= 16'hFFFF;
rommem[18474] <= 16'hFFFF;
rommem[18475] <= 16'hFFFF;
rommem[18476] <= 16'hFFFF;
rommem[18477] <= 16'hFFFF;
rommem[18478] <= 16'hFFFF;
rommem[18479] <= 16'hFFFF;
rommem[18480] <= 16'hFFFF;
rommem[18481] <= 16'hFFFF;
rommem[18482] <= 16'hFFFF;
rommem[18483] <= 16'hFFFF;
rommem[18484] <= 16'hFFFF;
rommem[18485] <= 16'hFFFF;
rommem[18486] <= 16'hFFFF;
rommem[18487] <= 16'hFFFF;
rommem[18488] <= 16'hFFFF;
rommem[18489] <= 16'hFFFF;
rommem[18490] <= 16'hFFFF;
rommem[18491] <= 16'hFFFF;
rommem[18492] <= 16'hFFFF;
rommem[18493] <= 16'hFFFF;
rommem[18494] <= 16'hFFFF;
rommem[18495] <= 16'hFFFF;
rommem[18496] <= 16'hFFFF;
rommem[18497] <= 16'hFFFF;
rommem[18498] <= 16'hFFFF;
rommem[18499] <= 16'hFFFF;
rommem[18500] <= 16'hFFFF;
rommem[18501] <= 16'hFFFF;
rommem[18502] <= 16'hFFFF;
rommem[18503] <= 16'hFFFF;
rommem[18504] <= 16'hFFFF;
rommem[18505] <= 16'hFFFF;
rommem[18506] <= 16'hFFFF;
rommem[18507] <= 16'hFFFF;
rommem[18508] <= 16'hFFFF;
rommem[18509] <= 16'hFFFF;
rommem[18510] <= 16'hFFFF;
rommem[18511] <= 16'hFFFF;
rommem[18512] <= 16'hFFFF;
rommem[18513] <= 16'hFFFF;
rommem[18514] <= 16'hFFFF;
rommem[18515] <= 16'hFFFF;
rommem[18516] <= 16'hFFFF;
rommem[18517] <= 16'hFFFF;
rommem[18518] <= 16'hFFFF;
rommem[18519] <= 16'hFFFF;
rommem[18520] <= 16'hFFFF;
rommem[18521] <= 16'hFFFF;
rommem[18522] <= 16'hFFFF;
rommem[18523] <= 16'hFFFF;
rommem[18524] <= 16'hFFFF;
rommem[18525] <= 16'hFFFF;
rommem[18526] <= 16'hFFFF;
rommem[18527] <= 16'hFFFF;
rommem[18528] <= 16'hFFFF;
rommem[18529] <= 16'hFFFF;
rommem[18530] <= 16'hFFFF;
rommem[18531] <= 16'hFFFF;
rommem[18532] <= 16'hFFFF;
rommem[18533] <= 16'hFFFF;
rommem[18534] <= 16'hFFFF;
rommem[18535] <= 16'hFFFF;
rommem[18536] <= 16'hFFFF;
rommem[18537] <= 16'hFFFF;
rommem[18538] <= 16'hFFFF;
rommem[18539] <= 16'hFFFF;
rommem[18540] <= 16'hFFFF;
rommem[18541] <= 16'hFFFF;
rommem[18542] <= 16'hFFFF;
rommem[18543] <= 16'hFFFF;
rommem[18544] <= 16'hFFFF;
rommem[18545] <= 16'hFFFF;
rommem[18546] <= 16'hFFFF;
rommem[18547] <= 16'hFFFF;
rommem[18548] <= 16'hFFFF;
rommem[18549] <= 16'hFFFF;
rommem[18550] <= 16'hFFFF;
rommem[18551] <= 16'hFFFF;
rommem[18552] <= 16'hFFFF;
rommem[18553] <= 16'hFFFF;
rommem[18554] <= 16'hFFFF;
rommem[18555] <= 16'hFFFF;
rommem[18556] <= 16'hFFFF;
rommem[18557] <= 16'hFFFF;
rommem[18558] <= 16'hFFFF;
rommem[18559] <= 16'hFFFF;
rommem[18560] <= 16'hFFFF;
rommem[18561] <= 16'hFFFF;
rommem[18562] <= 16'hFFFF;
rommem[18563] <= 16'hFFFF;
rommem[18564] <= 16'hFFFF;
rommem[18565] <= 16'hFFFF;
rommem[18566] <= 16'hFFFF;
rommem[18567] <= 16'hFFFF;
rommem[18568] <= 16'hFFFF;
rommem[18569] <= 16'hFFFF;
rommem[18570] <= 16'hFFFF;
rommem[18571] <= 16'hFFFF;
rommem[18572] <= 16'hFFFF;
rommem[18573] <= 16'hFFFF;
rommem[18574] <= 16'hFFFF;
rommem[18575] <= 16'hFFFF;
rommem[18576] <= 16'hFFFF;
rommem[18577] <= 16'hFFFF;
rommem[18578] <= 16'hFFFF;
rommem[18579] <= 16'hFFFF;
rommem[18580] <= 16'hFFFF;
rommem[18581] <= 16'hFFFF;
rommem[18582] <= 16'hFFFF;
rommem[18583] <= 16'hFFFF;
rommem[18584] <= 16'hFFFF;
rommem[18585] <= 16'hFFFF;
rommem[18586] <= 16'hFFFF;
rommem[18587] <= 16'hFFFF;
rommem[18588] <= 16'hFFFF;
rommem[18589] <= 16'hFFFF;
rommem[18590] <= 16'hFFFF;
rommem[18591] <= 16'hFFFF;
rommem[18592] <= 16'hFFFF;
rommem[18593] <= 16'hFFFF;
rommem[18594] <= 16'hFFFF;
rommem[18595] <= 16'hFFFF;
rommem[18596] <= 16'hFFFF;
rommem[18597] <= 16'hFFFF;
rommem[18598] <= 16'hFFFF;
rommem[18599] <= 16'hFFFF;
rommem[18600] <= 16'hFFFF;
rommem[18601] <= 16'hFFFF;
rommem[18602] <= 16'hFFFF;
rommem[18603] <= 16'hFFFF;
rommem[18604] <= 16'hFFFF;
rommem[18605] <= 16'hFFFF;
rommem[18606] <= 16'hFFFF;
rommem[18607] <= 16'hFFFF;
rommem[18608] <= 16'hFFFF;
rommem[18609] <= 16'hFFFF;
rommem[18610] <= 16'hFFFF;
rommem[18611] <= 16'hFFFF;
rommem[18612] <= 16'hFFFF;
rommem[18613] <= 16'hFFFF;
rommem[18614] <= 16'hFFFF;
rommem[18615] <= 16'hFFFF;
rommem[18616] <= 16'hFFFF;
rommem[18617] <= 16'hFFFF;
rommem[18618] <= 16'hFFFF;
rommem[18619] <= 16'hFFFF;
rommem[18620] <= 16'hFFFF;
rommem[18621] <= 16'hFFFF;
rommem[18622] <= 16'hFFFF;
rommem[18623] <= 16'hFFFF;
rommem[18624] <= 16'hFFFF;
rommem[18625] <= 16'hFFFF;
rommem[18626] <= 16'hFFFF;
rommem[18627] <= 16'hFFFF;
rommem[18628] <= 16'hFFFF;
rommem[18629] <= 16'hFFFF;
rommem[18630] <= 16'hFFFF;
rommem[18631] <= 16'hFFFF;
rommem[18632] <= 16'hFFFF;
rommem[18633] <= 16'hFFFF;
rommem[18634] <= 16'hFFFF;
rommem[18635] <= 16'hFFFF;
rommem[18636] <= 16'hFFFF;
rommem[18637] <= 16'hFFFF;
rommem[18638] <= 16'hFFFF;
rommem[18639] <= 16'hFFFF;
rommem[18640] <= 16'hFFFF;
rommem[18641] <= 16'hFFFF;
rommem[18642] <= 16'hFFFF;
rommem[18643] <= 16'hFFFF;
rommem[18644] <= 16'hFFFF;
rommem[18645] <= 16'hFFFF;
rommem[18646] <= 16'hFFFF;
rommem[18647] <= 16'hFFFF;
rommem[18648] <= 16'hFFFF;
rommem[18649] <= 16'hFFFF;
rommem[18650] <= 16'hFFFF;
rommem[18651] <= 16'hFFFF;
rommem[18652] <= 16'hFFFF;
rommem[18653] <= 16'hFFFF;
rommem[18654] <= 16'hFFFF;
rommem[18655] <= 16'hFFFF;
rommem[18656] <= 16'hFFFF;
rommem[18657] <= 16'hFFFF;
rommem[18658] <= 16'hFFFF;
rommem[18659] <= 16'hFFFF;
rommem[18660] <= 16'hFFFF;
rommem[18661] <= 16'hFFFF;
rommem[18662] <= 16'hFFFF;
rommem[18663] <= 16'hFFFF;
rommem[18664] <= 16'hFFFF;
rommem[18665] <= 16'hFFFF;
rommem[18666] <= 16'hFFFF;
rommem[18667] <= 16'hFFFF;
rommem[18668] <= 16'hFFFF;
rommem[18669] <= 16'hFFFF;
rommem[18670] <= 16'hFFFF;
rommem[18671] <= 16'hFFFF;
rommem[18672] <= 16'hFFFF;
rommem[18673] <= 16'hFFFF;
rommem[18674] <= 16'hFFFF;
rommem[18675] <= 16'hFFFF;
rommem[18676] <= 16'hFFFF;
rommem[18677] <= 16'hFFFF;
rommem[18678] <= 16'hFFFF;
rommem[18679] <= 16'hFFFF;
rommem[18680] <= 16'hFFFF;
rommem[18681] <= 16'hFFFF;
rommem[18682] <= 16'hFFFF;
rommem[18683] <= 16'hFFFF;
rommem[18684] <= 16'hFFFF;
rommem[18685] <= 16'hFFFF;
rommem[18686] <= 16'hFFFF;
rommem[18687] <= 16'hFFFF;
rommem[18688] <= 16'hFFFF;
rommem[18689] <= 16'hFFFF;
rommem[18690] <= 16'hFFFF;
rommem[18691] <= 16'hFFFF;
rommem[18692] <= 16'hFFFF;
rommem[18693] <= 16'hFFFF;
rommem[18694] <= 16'hFFFF;
rommem[18695] <= 16'hFFFF;
rommem[18696] <= 16'hFFFF;
rommem[18697] <= 16'hFFFF;
rommem[18698] <= 16'hFFFF;
rommem[18699] <= 16'hFFFF;
rommem[18700] <= 16'hFFFF;
rommem[18701] <= 16'hFFFF;
rommem[18702] <= 16'hFFFF;
rommem[18703] <= 16'hFFFF;
rommem[18704] <= 16'hFFFF;
rommem[18705] <= 16'hFFFF;
rommem[18706] <= 16'hFFFF;
rommem[18707] <= 16'hFFFF;
rommem[18708] <= 16'hFFFF;
rommem[18709] <= 16'hFFFF;
rommem[18710] <= 16'hFFFF;
rommem[18711] <= 16'hFFFF;
rommem[18712] <= 16'hFFFF;
rommem[18713] <= 16'hFFFF;
rommem[18714] <= 16'hFFFF;
rommem[18715] <= 16'hFFFF;
rommem[18716] <= 16'hFFFF;
rommem[18717] <= 16'hFFFF;
rommem[18718] <= 16'hFFFF;
rommem[18719] <= 16'hFFFF;
rommem[18720] <= 16'hFFFF;
rommem[18721] <= 16'hFFFF;
rommem[18722] <= 16'hFFFF;
rommem[18723] <= 16'hFFFF;
rommem[18724] <= 16'hFFFF;
rommem[18725] <= 16'hFFFF;
rommem[18726] <= 16'hFFFF;
rommem[18727] <= 16'hFFFF;
rommem[18728] <= 16'hFFFF;
rommem[18729] <= 16'hFFFF;
rommem[18730] <= 16'hFFFF;
rommem[18731] <= 16'hFFFF;
rommem[18732] <= 16'hFFFF;
rommem[18733] <= 16'hFFFF;
rommem[18734] <= 16'hFFFF;
rommem[18735] <= 16'hFFFF;
rommem[18736] <= 16'hFFFF;
rommem[18737] <= 16'hFFFF;
rommem[18738] <= 16'hFFFF;
rommem[18739] <= 16'hFFFF;
rommem[18740] <= 16'hFFFF;
rommem[18741] <= 16'hFFFF;
rommem[18742] <= 16'hFFFF;
rommem[18743] <= 16'hFFFF;
rommem[18744] <= 16'hFFFF;
rommem[18745] <= 16'hFFFF;
rommem[18746] <= 16'hFFFF;
rommem[18747] <= 16'hFFFF;
rommem[18748] <= 16'hFFFF;
rommem[18749] <= 16'hFFFF;
rommem[18750] <= 16'hFFFF;
rommem[18751] <= 16'hFFFF;
rommem[18752] <= 16'hFFFF;
rommem[18753] <= 16'hFFFF;
rommem[18754] <= 16'hFFFF;
rommem[18755] <= 16'hFFFF;
rommem[18756] <= 16'hFFFF;
rommem[18757] <= 16'hFFFF;
rommem[18758] <= 16'hFFFF;
rommem[18759] <= 16'hFFFF;
rommem[18760] <= 16'hFFFF;
rommem[18761] <= 16'hFFFF;
rommem[18762] <= 16'hFFFF;
rommem[18763] <= 16'hFFFF;
rommem[18764] <= 16'hFFFF;
rommem[18765] <= 16'hFFFF;
rommem[18766] <= 16'hFFFF;
rommem[18767] <= 16'hFFFF;
rommem[18768] <= 16'hFFFF;
rommem[18769] <= 16'hFFFF;
rommem[18770] <= 16'hFFFF;
rommem[18771] <= 16'hFFFF;
rommem[18772] <= 16'hFFFF;
rommem[18773] <= 16'hFFFF;
rommem[18774] <= 16'hFFFF;
rommem[18775] <= 16'hFFFF;
rommem[18776] <= 16'hFFFF;
rommem[18777] <= 16'hFFFF;
rommem[18778] <= 16'hFFFF;
rommem[18779] <= 16'hFFFF;
rommem[18780] <= 16'hFFFF;
rommem[18781] <= 16'hFFFF;
rommem[18782] <= 16'hFFFF;
rommem[18783] <= 16'hFFFF;
rommem[18784] <= 16'hFFFF;
rommem[18785] <= 16'hFFFF;
rommem[18786] <= 16'hFFFF;
rommem[18787] <= 16'hFFFF;
rommem[18788] <= 16'hFFFF;
rommem[18789] <= 16'hFFFF;
rommem[18790] <= 16'hFFFF;
rommem[18791] <= 16'hFFFF;
rommem[18792] <= 16'hFFFF;
rommem[18793] <= 16'hFFFF;
rommem[18794] <= 16'hFFFF;
rommem[18795] <= 16'hFFFF;
rommem[18796] <= 16'hFFFF;
rommem[18797] <= 16'hFFFF;
rommem[18798] <= 16'hFFFF;
rommem[18799] <= 16'hFFFF;
rommem[18800] <= 16'hFFFF;
rommem[18801] <= 16'hFFFF;
rommem[18802] <= 16'hFFFF;
rommem[18803] <= 16'hFFFF;
rommem[18804] <= 16'hFFFF;
rommem[18805] <= 16'hFFFF;
rommem[18806] <= 16'hFFFF;
rommem[18807] <= 16'hFFFF;
rommem[18808] <= 16'hFFFF;
rommem[18809] <= 16'hFFFF;
rommem[18810] <= 16'hFFFF;
rommem[18811] <= 16'hFFFF;
rommem[18812] <= 16'hFFFF;
rommem[18813] <= 16'hFFFF;
rommem[18814] <= 16'hFFFF;
rommem[18815] <= 16'hFFFF;
rommem[18816] <= 16'hFFFF;
rommem[18817] <= 16'hFFFF;
rommem[18818] <= 16'hFFFF;
rommem[18819] <= 16'hFFFF;
rommem[18820] <= 16'hFFFF;
rommem[18821] <= 16'hFFFF;
rommem[18822] <= 16'hFFFF;
rommem[18823] <= 16'hFFFF;
rommem[18824] <= 16'hFFFF;
rommem[18825] <= 16'hFFFF;
rommem[18826] <= 16'hFFFF;
rommem[18827] <= 16'hFFFF;
rommem[18828] <= 16'hFFFF;
rommem[18829] <= 16'hFFFF;
rommem[18830] <= 16'hFFFF;
rommem[18831] <= 16'hFFFF;
rommem[18832] <= 16'hFFFF;
rommem[18833] <= 16'hFFFF;
rommem[18834] <= 16'hFFFF;
rommem[18835] <= 16'hFFFF;
rommem[18836] <= 16'hFFFF;
rommem[18837] <= 16'hFFFF;
rommem[18838] <= 16'hFFFF;
rommem[18839] <= 16'hFFFF;
rommem[18840] <= 16'hFFFF;
rommem[18841] <= 16'hFFFF;
rommem[18842] <= 16'hFFFF;
rommem[18843] <= 16'hFFFF;
rommem[18844] <= 16'hFFFF;
rommem[18845] <= 16'hFFFF;
rommem[18846] <= 16'hFFFF;
rommem[18847] <= 16'hFFFF;
rommem[18848] <= 16'hFFFF;
rommem[18849] <= 16'hFFFF;
rommem[18850] <= 16'hFFFF;
rommem[18851] <= 16'hFFFF;
rommem[18852] <= 16'hFFFF;
rommem[18853] <= 16'hFFFF;
rommem[18854] <= 16'hFFFF;
rommem[18855] <= 16'hFFFF;
rommem[18856] <= 16'hFFFF;
rommem[18857] <= 16'hFFFF;
rommem[18858] <= 16'hFFFF;
rommem[18859] <= 16'hFFFF;
rommem[18860] <= 16'hFFFF;
rommem[18861] <= 16'hFFFF;
rommem[18862] <= 16'hFFFF;
rommem[18863] <= 16'hFFFF;
rommem[18864] <= 16'hFFFF;
rommem[18865] <= 16'hFFFF;
rommem[18866] <= 16'hFFFF;
rommem[18867] <= 16'hFFFF;
rommem[18868] <= 16'hFFFF;
rommem[18869] <= 16'hFFFF;
rommem[18870] <= 16'hFFFF;
rommem[18871] <= 16'hFFFF;
rommem[18872] <= 16'hFFFF;
rommem[18873] <= 16'hFFFF;
rommem[18874] <= 16'hFFFF;
rommem[18875] <= 16'hFFFF;
rommem[18876] <= 16'hFFFF;
rommem[18877] <= 16'hFFFF;
rommem[18878] <= 16'hFFFF;
rommem[18879] <= 16'hFFFF;
rommem[18880] <= 16'hFFFF;
rommem[18881] <= 16'hFFFF;
rommem[18882] <= 16'hFFFF;
rommem[18883] <= 16'hFFFF;
rommem[18884] <= 16'hFFFF;
rommem[18885] <= 16'hFFFF;
rommem[18886] <= 16'hFFFF;
rommem[18887] <= 16'hFFFF;
rommem[18888] <= 16'hFFFF;
rommem[18889] <= 16'hFFFF;
rommem[18890] <= 16'hFFFF;
rommem[18891] <= 16'hFFFF;
rommem[18892] <= 16'hFFFF;
rommem[18893] <= 16'hFFFF;
rommem[18894] <= 16'hFFFF;
rommem[18895] <= 16'hFFFF;
rommem[18896] <= 16'hFFFF;
rommem[18897] <= 16'hFFFF;
rommem[18898] <= 16'hFFFF;
rommem[18899] <= 16'hFFFF;
rommem[18900] <= 16'hFFFF;
rommem[18901] <= 16'hFFFF;
rommem[18902] <= 16'hFFFF;
rommem[18903] <= 16'hFFFF;
rommem[18904] <= 16'hFFFF;
rommem[18905] <= 16'hFFFF;
rommem[18906] <= 16'hFFFF;
rommem[18907] <= 16'hFFFF;
rommem[18908] <= 16'hFFFF;
rommem[18909] <= 16'hFFFF;
rommem[18910] <= 16'hFFFF;
rommem[18911] <= 16'hFFFF;
rommem[18912] <= 16'hFFFF;
rommem[18913] <= 16'hFFFF;
rommem[18914] <= 16'hFFFF;
rommem[18915] <= 16'hFFFF;
rommem[18916] <= 16'hFFFF;
rommem[18917] <= 16'hFFFF;
rommem[18918] <= 16'hFFFF;
rommem[18919] <= 16'hFFFF;
rommem[18920] <= 16'hFFFF;
rommem[18921] <= 16'hFFFF;
rommem[18922] <= 16'hFFFF;
rommem[18923] <= 16'hFFFF;
rommem[18924] <= 16'hFFFF;
rommem[18925] <= 16'hFFFF;
rommem[18926] <= 16'hFFFF;
rommem[18927] <= 16'hFFFF;
rommem[18928] <= 16'hFFFF;
rommem[18929] <= 16'hFFFF;
rommem[18930] <= 16'hFFFF;
rommem[18931] <= 16'hFFFF;
rommem[18932] <= 16'hFFFF;
rommem[18933] <= 16'hFFFF;
rommem[18934] <= 16'hFFFF;
rommem[18935] <= 16'hFFFF;
rommem[18936] <= 16'hFFFF;
rommem[18937] <= 16'hFFFF;
rommem[18938] <= 16'hFFFF;
rommem[18939] <= 16'hFFFF;
rommem[18940] <= 16'hFFFF;
rommem[18941] <= 16'hFFFF;
rommem[18942] <= 16'hFFFF;
rommem[18943] <= 16'hFFFF;
rommem[18944] <= 16'hFFFF;
rommem[18945] <= 16'hFFFF;
rommem[18946] <= 16'hFFFF;
rommem[18947] <= 16'hFFFF;
rommem[18948] <= 16'hFFFF;
rommem[18949] <= 16'hFFFF;
rommem[18950] <= 16'hFFFF;
rommem[18951] <= 16'hFFFF;
rommem[18952] <= 16'hFFFF;
rommem[18953] <= 16'hFFFF;
rommem[18954] <= 16'hFFFF;
rommem[18955] <= 16'hFFFF;
rommem[18956] <= 16'hFFFF;
rommem[18957] <= 16'hFFFF;
rommem[18958] <= 16'hFFFF;
rommem[18959] <= 16'hFFFF;
rommem[18960] <= 16'hFFFF;
rommem[18961] <= 16'hFFFF;
rommem[18962] <= 16'hFFFF;
rommem[18963] <= 16'hFFFF;
rommem[18964] <= 16'hFFFF;
rommem[18965] <= 16'hFFFF;
rommem[18966] <= 16'hFFFF;
rommem[18967] <= 16'hFFFF;
rommem[18968] <= 16'hFFFF;
rommem[18969] <= 16'hFFFF;
rommem[18970] <= 16'hFFFF;
rommem[18971] <= 16'hFFFF;
rommem[18972] <= 16'hFFFF;
rommem[18973] <= 16'hFFFF;
rommem[18974] <= 16'hFFFF;
rommem[18975] <= 16'hFFFF;
rommem[18976] <= 16'hFFFF;
rommem[18977] <= 16'hFFFF;
rommem[18978] <= 16'hFFFF;
rommem[18979] <= 16'hFFFF;
rommem[18980] <= 16'hFFFF;
rommem[18981] <= 16'hFFFF;
rommem[18982] <= 16'hFFFF;
rommem[18983] <= 16'hFFFF;
rommem[18984] <= 16'hFFFF;
rommem[18985] <= 16'hFFFF;
rommem[18986] <= 16'hFFFF;
rommem[18987] <= 16'hFFFF;
rommem[18988] <= 16'hFFFF;
rommem[18989] <= 16'hFFFF;
rommem[18990] <= 16'hFFFF;
rommem[18991] <= 16'hFFFF;
rommem[18992] <= 16'hFFFF;
rommem[18993] <= 16'hFFFF;
rommem[18994] <= 16'hFFFF;
rommem[18995] <= 16'hFFFF;
rommem[18996] <= 16'hFFFF;
rommem[18997] <= 16'hFFFF;
rommem[18998] <= 16'hFFFF;
rommem[18999] <= 16'hFFFF;
rommem[19000] <= 16'hFFFF;
rommem[19001] <= 16'hFFFF;
rommem[19002] <= 16'hFFFF;
rommem[19003] <= 16'hFFFF;
rommem[19004] <= 16'hFFFF;
rommem[19005] <= 16'hFFFF;
rommem[19006] <= 16'hFFFF;
rommem[19007] <= 16'hFFFF;
rommem[19008] <= 16'hFFFF;
rommem[19009] <= 16'hFFFF;
rommem[19010] <= 16'hFFFF;
rommem[19011] <= 16'hFFFF;
rommem[19012] <= 16'hFFFF;
rommem[19013] <= 16'hFFFF;
rommem[19014] <= 16'hFFFF;
rommem[19015] <= 16'hFFFF;
rommem[19016] <= 16'hFFFF;
rommem[19017] <= 16'hFFFF;
rommem[19018] <= 16'hFFFF;
rommem[19019] <= 16'hFFFF;
rommem[19020] <= 16'hFFFF;
rommem[19021] <= 16'hFFFF;
rommem[19022] <= 16'hFFFF;
rommem[19023] <= 16'hFFFF;
rommem[19024] <= 16'hFFFF;
rommem[19025] <= 16'hFFFF;
rommem[19026] <= 16'hFFFF;
rommem[19027] <= 16'hFFFF;
rommem[19028] <= 16'hFFFF;
rommem[19029] <= 16'hFFFF;
rommem[19030] <= 16'hFFFF;
rommem[19031] <= 16'hFFFF;
rommem[19032] <= 16'hFFFF;
rommem[19033] <= 16'hFFFF;
rommem[19034] <= 16'hFFFF;
rommem[19035] <= 16'hFFFF;
rommem[19036] <= 16'hFFFF;
rommem[19037] <= 16'hFFFF;
rommem[19038] <= 16'hFFFF;
rommem[19039] <= 16'hFFFF;
rommem[19040] <= 16'hFFFF;
rommem[19041] <= 16'hFFFF;
rommem[19042] <= 16'hFFFF;
rommem[19043] <= 16'hFFFF;
rommem[19044] <= 16'hFFFF;
rommem[19045] <= 16'hFFFF;
rommem[19046] <= 16'hFFFF;
rommem[19047] <= 16'hFFFF;
rommem[19048] <= 16'hFFFF;
rommem[19049] <= 16'hFFFF;
rommem[19050] <= 16'hFFFF;
rommem[19051] <= 16'hFFFF;
rommem[19052] <= 16'hFFFF;
rommem[19053] <= 16'hFFFF;
rommem[19054] <= 16'hFFFF;
rommem[19055] <= 16'hFFFF;
rommem[19056] <= 16'hFFFF;
rommem[19057] <= 16'hFFFF;
rommem[19058] <= 16'hFFFF;
rommem[19059] <= 16'hFFFF;
rommem[19060] <= 16'hFFFF;
rommem[19061] <= 16'hFFFF;
rommem[19062] <= 16'hFFFF;
rommem[19063] <= 16'hFFFF;
rommem[19064] <= 16'hFFFF;
rommem[19065] <= 16'hFFFF;
rommem[19066] <= 16'hFFFF;
rommem[19067] <= 16'hFFFF;
rommem[19068] <= 16'hFFFF;
rommem[19069] <= 16'hFFFF;
rommem[19070] <= 16'hFFFF;
rommem[19071] <= 16'hFFFF;
rommem[19072] <= 16'hFFFF;
rommem[19073] <= 16'hFFFF;
rommem[19074] <= 16'hFFFF;
rommem[19075] <= 16'hFFFF;
rommem[19076] <= 16'hFFFF;
rommem[19077] <= 16'hFFFF;
rommem[19078] <= 16'hFFFF;
rommem[19079] <= 16'hFFFF;
rommem[19080] <= 16'hFFFF;
rommem[19081] <= 16'hFFFF;
rommem[19082] <= 16'hFFFF;
rommem[19083] <= 16'hFFFF;
rommem[19084] <= 16'hFFFF;
rommem[19085] <= 16'hFFFF;
rommem[19086] <= 16'hFFFF;
rommem[19087] <= 16'hFFFF;
rommem[19088] <= 16'hFFFF;
rommem[19089] <= 16'hFFFF;
rommem[19090] <= 16'hFFFF;
rommem[19091] <= 16'hFFFF;
rommem[19092] <= 16'hFFFF;
rommem[19093] <= 16'hFFFF;
rommem[19094] <= 16'hFFFF;
rommem[19095] <= 16'hFFFF;
rommem[19096] <= 16'hFFFF;
rommem[19097] <= 16'hFFFF;
rommem[19098] <= 16'hFFFF;
rommem[19099] <= 16'hFFFF;
rommem[19100] <= 16'hFFFF;
rommem[19101] <= 16'hFFFF;
rommem[19102] <= 16'hFFFF;
rommem[19103] <= 16'hFFFF;
rommem[19104] <= 16'hFFFF;
rommem[19105] <= 16'hFFFF;
rommem[19106] <= 16'hFFFF;
rommem[19107] <= 16'hFFFF;
rommem[19108] <= 16'hFFFF;
rommem[19109] <= 16'hFFFF;
rommem[19110] <= 16'hFFFF;
rommem[19111] <= 16'hFFFF;
rommem[19112] <= 16'hFFFF;
rommem[19113] <= 16'hFFFF;
rommem[19114] <= 16'hFFFF;
rommem[19115] <= 16'hFFFF;
rommem[19116] <= 16'hFFFF;
rommem[19117] <= 16'hFFFF;
rommem[19118] <= 16'hFFFF;
rommem[19119] <= 16'hFFFF;
rommem[19120] <= 16'hFFFF;
rommem[19121] <= 16'hFFFF;
rommem[19122] <= 16'hFFFF;
rommem[19123] <= 16'hFFFF;
rommem[19124] <= 16'hFFFF;
rommem[19125] <= 16'hFFFF;
rommem[19126] <= 16'hFFFF;
rommem[19127] <= 16'hFFFF;
rommem[19128] <= 16'hFFFF;
rommem[19129] <= 16'hFFFF;
rommem[19130] <= 16'hFFFF;
rommem[19131] <= 16'hFFFF;
rommem[19132] <= 16'hFFFF;
rommem[19133] <= 16'hFFFF;
rommem[19134] <= 16'hFFFF;
rommem[19135] <= 16'hFFFF;
rommem[19136] <= 16'hFFFF;
rommem[19137] <= 16'hFFFF;
rommem[19138] <= 16'hFFFF;
rommem[19139] <= 16'hFFFF;
rommem[19140] <= 16'hFFFF;
rommem[19141] <= 16'hFFFF;
rommem[19142] <= 16'hFFFF;
rommem[19143] <= 16'hFFFF;
rommem[19144] <= 16'hFFFF;
rommem[19145] <= 16'hFFFF;
rommem[19146] <= 16'hFFFF;
rommem[19147] <= 16'hFFFF;
rommem[19148] <= 16'hFFFF;
rommem[19149] <= 16'hFFFF;
rommem[19150] <= 16'hFFFF;
rommem[19151] <= 16'hFFFF;
rommem[19152] <= 16'hFFFF;
rommem[19153] <= 16'hFFFF;
rommem[19154] <= 16'hFFFF;
rommem[19155] <= 16'hFFFF;
rommem[19156] <= 16'hFFFF;
rommem[19157] <= 16'hFFFF;
rommem[19158] <= 16'hFFFF;
rommem[19159] <= 16'hFFFF;
rommem[19160] <= 16'hFFFF;
rommem[19161] <= 16'hFFFF;
rommem[19162] <= 16'hFFFF;
rommem[19163] <= 16'hFFFF;
rommem[19164] <= 16'hFFFF;
rommem[19165] <= 16'hFFFF;
rommem[19166] <= 16'hFFFF;
rommem[19167] <= 16'hFFFF;
rommem[19168] <= 16'hFFFF;
rommem[19169] <= 16'hFFFF;
rommem[19170] <= 16'hFFFF;
rommem[19171] <= 16'hFFFF;
rommem[19172] <= 16'hFFFF;
rommem[19173] <= 16'hFFFF;
rommem[19174] <= 16'hFFFF;
rommem[19175] <= 16'hFFFF;
rommem[19176] <= 16'hFFFF;
rommem[19177] <= 16'hFFFF;
rommem[19178] <= 16'hFFFF;
rommem[19179] <= 16'hFFFF;
rommem[19180] <= 16'hFFFF;
rommem[19181] <= 16'hFFFF;
rommem[19182] <= 16'hFFFF;
rommem[19183] <= 16'hFFFF;
rommem[19184] <= 16'hFFFF;
rommem[19185] <= 16'hFFFF;
rommem[19186] <= 16'hFFFF;
rommem[19187] <= 16'hFFFF;
rommem[19188] <= 16'hFFFF;
rommem[19189] <= 16'hFFFF;
rommem[19190] <= 16'hFFFF;
rommem[19191] <= 16'hFFFF;
rommem[19192] <= 16'hFFFF;
rommem[19193] <= 16'hFFFF;
rommem[19194] <= 16'hFFFF;
rommem[19195] <= 16'hFFFF;
rommem[19196] <= 16'hFFFF;
rommem[19197] <= 16'hFFFF;
rommem[19198] <= 16'hFFFF;
rommem[19199] <= 16'hFFFF;
rommem[19200] <= 16'hFFFF;
rommem[19201] <= 16'hFFFF;
rommem[19202] <= 16'hFFFF;
rommem[19203] <= 16'hFFFF;
rommem[19204] <= 16'hFFFF;
rommem[19205] <= 16'hFFFF;
rommem[19206] <= 16'hFFFF;
rommem[19207] <= 16'hFFFF;
rommem[19208] <= 16'hFFFF;
rommem[19209] <= 16'hFFFF;
rommem[19210] <= 16'hFFFF;
rommem[19211] <= 16'hFFFF;
rommem[19212] <= 16'hFFFF;
rommem[19213] <= 16'hFFFF;
rommem[19214] <= 16'hFFFF;
rommem[19215] <= 16'hFFFF;
rommem[19216] <= 16'hFFFF;
rommem[19217] <= 16'hFFFF;
rommem[19218] <= 16'hFFFF;
rommem[19219] <= 16'hFFFF;
rommem[19220] <= 16'hFFFF;
rommem[19221] <= 16'hFFFF;
rommem[19222] <= 16'hFFFF;
rommem[19223] <= 16'hFFFF;
rommem[19224] <= 16'hFFFF;
rommem[19225] <= 16'hFFFF;
rommem[19226] <= 16'hFFFF;
rommem[19227] <= 16'hFFFF;
rommem[19228] <= 16'hFFFF;
rommem[19229] <= 16'hFFFF;
rommem[19230] <= 16'hFFFF;
rommem[19231] <= 16'hFFFF;
rommem[19232] <= 16'hFFFF;
rommem[19233] <= 16'hFFFF;
rommem[19234] <= 16'hFFFF;
rommem[19235] <= 16'hFFFF;
rommem[19236] <= 16'hFFFF;
rommem[19237] <= 16'hFFFF;
rommem[19238] <= 16'hFFFF;
rommem[19239] <= 16'hFFFF;
rommem[19240] <= 16'hFFFF;
rommem[19241] <= 16'hFFFF;
rommem[19242] <= 16'hFFFF;
rommem[19243] <= 16'hFFFF;
rommem[19244] <= 16'hFFFF;
rommem[19245] <= 16'hFFFF;
rommem[19246] <= 16'hFFFF;
rommem[19247] <= 16'hFFFF;
rommem[19248] <= 16'hFFFF;
rommem[19249] <= 16'hFFFF;
rommem[19250] <= 16'hFFFF;
rommem[19251] <= 16'hFFFF;
rommem[19252] <= 16'hFFFF;
rommem[19253] <= 16'hFFFF;
rommem[19254] <= 16'hFFFF;
rommem[19255] <= 16'hFFFF;
rommem[19256] <= 16'hFFFF;
rommem[19257] <= 16'hFFFF;
rommem[19258] <= 16'hFFFF;
rommem[19259] <= 16'hFFFF;
rommem[19260] <= 16'hFFFF;
rommem[19261] <= 16'hFFFF;
rommem[19262] <= 16'hFFFF;
rommem[19263] <= 16'hFFFF;
rommem[19264] <= 16'hFFFF;
rommem[19265] <= 16'hFFFF;
rommem[19266] <= 16'hFFFF;
rommem[19267] <= 16'hFFFF;
rommem[19268] <= 16'hFFFF;
rommem[19269] <= 16'hFFFF;
rommem[19270] <= 16'hFFFF;
rommem[19271] <= 16'hFFFF;
rommem[19272] <= 16'hFFFF;
rommem[19273] <= 16'hFFFF;
rommem[19274] <= 16'hFFFF;
rommem[19275] <= 16'hFFFF;
rommem[19276] <= 16'hFFFF;
rommem[19277] <= 16'hFFFF;
rommem[19278] <= 16'hFFFF;
rommem[19279] <= 16'hFFFF;
rommem[19280] <= 16'hFFFF;
rommem[19281] <= 16'hFFFF;
rommem[19282] <= 16'hFFFF;
rommem[19283] <= 16'hFFFF;
rommem[19284] <= 16'hFFFF;
rommem[19285] <= 16'hFFFF;
rommem[19286] <= 16'hFFFF;
rommem[19287] <= 16'hFFFF;
rommem[19288] <= 16'hFFFF;
rommem[19289] <= 16'hFFFF;
rommem[19290] <= 16'hFFFF;
rommem[19291] <= 16'hFFFF;
rommem[19292] <= 16'hFFFF;
rommem[19293] <= 16'hFFFF;
rommem[19294] <= 16'hFFFF;
rommem[19295] <= 16'hFFFF;
rommem[19296] <= 16'hFFFF;
rommem[19297] <= 16'hFFFF;
rommem[19298] <= 16'hFFFF;
rommem[19299] <= 16'hFFFF;
rommem[19300] <= 16'hFFFF;
rommem[19301] <= 16'hFFFF;
rommem[19302] <= 16'hFFFF;
rommem[19303] <= 16'hFFFF;
rommem[19304] <= 16'hFFFF;
rommem[19305] <= 16'hFFFF;
rommem[19306] <= 16'hFFFF;
rommem[19307] <= 16'hFFFF;
rommem[19308] <= 16'hFFFF;
rommem[19309] <= 16'hFFFF;
rommem[19310] <= 16'hFFFF;
rommem[19311] <= 16'hFFFF;
rommem[19312] <= 16'hFFFF;
rommem[19313] <= 16'hFFFF;
rommem[19314] <= 16'hFFFF;
rommem[19315] <= 16'hFFFF;
rommem[19316] <= 16'hFFFF;
rommem[19317] <= 16'hFFFF;
rommem[19318] <= 16'hFFFF;
rommem[19319] <= 16'hFFFF;
rommem[19320] <= 16'hFFFF;
rommem[19321] <= 16'hFFFF;
rommem[19322] <= 16'hFFFF;
rommem[19323] <= 16'hFFFF;
rommem[19324] <= 16'hFFFF;
rommem[19325] <= 16'hFFFF;
rommem[19326] <= 16'hFFFF;
rommem[19327] <= 16'hFFFF;
rommem[19328] <= 16'hFFFF;
rommem[19329] <= 16'hFFFF;
rommem[19330] <= 16'hFFFF;
rommem[19331] <= 16'hFFFF;
rommem[19332] <= 16'hFFFF;
rommem[19333] <= 16'hFFFF;
rommem[19334] <= 16'hFFFF;
rommem[19335] <= 16'hFFFF;
rommem[19336] <= 16'hFFFF;
rommem[19337] <= 16'hFFFF;
rommem[19338] <= 16'hFFFF;
rommem[19339] <= 16'hFFFF;
rommem[19340] <= 16'hFFFF;
rommem[19341] <= 16'hFFFF;
rommem[19342] <= 16'hFFFF;
rommem[19343] <= 16'hFFFF;
rommem[19344] <= 16'hFFFF;
rommem[19345] <= 16'hFFFF;
rommem[19346] <= 16'hFFFF;
rommem[19347] <= 16'hFFFF;
rommem[19348] <= 16'hFFFF;
rommem[19349] <= 16'hFFFF;
rommem[19350] <= 16'hFFFF;
rommem[19351] <= 16'hFFFF;
rommem[19352] <= 16'hFFFF;
rommem[19353] <= 16'hFFFF;
rommem[19354] <= 16'hFFFF;
rommem[19355] <= 16'hFFFF;
rommem[19356] <= 16'hFFFF;
rommem[19357] <= 16'hFFFF;
rommem[19358] <= 16'hFFFF;
rommem[19359] <= 16'hFFFF;
rommem[19360] <= 16'hFFFF;
rommem[19361] <= 16'hFFFF;
rommem[19362] <= 16'hFFFF;
rommem[19363] <= 16'hFFFF;
rommem[19364] <= 16'hFFFF;
rommem[19365] <= 16'hFFFF;
rommem[19366] <= 16'hFFFF;
rommem[19367] <= 16'hFFFF;
rommem[19368] <= 16'hFFFF;
rommem[19369] <= 16'hFFFF;
rommem[19370] <= 16'hFFFF;
rommem[19371] <= 16'hFFFF;
rommem[19372] <= 16'hFFFF;
rommem[19373] <= 16'hFFFF;
rommem[19374] <= 16'hFFFF;
rommem[19375] <= 16'hFFFF;
rommem[19376] <= 16'hFFFF;
rommem[19377] <= 16'hFFFF;
rommem[19378] <= 16'hFFFF;
rommem[19379] <= 16'hFFFF;
rommem[19380] <= 16'hFFFF;
rommem[19381] <= 16'hFFFF;
rommem[19382] <= 16'hFFFF;
rommem[19383] <= 16'hFFFF;
rommem[19384] <= 16'hFFFF;
rommem[19385] <= 16'hFFFF;
rommem[19386] <= 16'hFFFF;
rommem[19387] <= 16'hFFFF;
rommem[19388] <= 16'hFFFF;
rommem[19389] <= 16'hFFFF;
rommem[19390] <= 16'hFFFF;
rommem[19391] <= 16'hFFFF;
rommem[19392] <= 16'hFFFF;
rommem[19393] <= 16'hFFFF;
rommem[19394] <= 16'hFFFF;
rommem[19395] <= 16'hFFFF;
rommem[19396] <= 16'hFFFF;
rommem[19397] <= 16'hFFFF;
rommem[19398] <= 16'hFFFF;
rommem[19399] <= 16'hFFFF;
rommem[19400] <= 16'hFFFF;
rommem[19401] <= 16'hFFFF;
rommem[19402] <= 16'hFFFF;
rommem[19403] <= 16'hFFFF;
rommem[19404] <= 16'hFFFF;
rommem[19405] <= 16'hFFFF;
rommem[19406] <= 16'hFFFF;
rommem[19407] <= 16'hFFFF;
rommem[19408] <= 16'hFFFF;
rommem[19409] <= 16'hFFFF;
rommem[19410] <= 16'hFFFF;
rommem[19411] <= 16'hFFFF;
rommem[19412] <= 16'hFFFF;
rommem[19413] <= 16'hFFFF;
rommem[19414] <= 16'hFFFF;
rommem[19415] <= 16'hFFFF;
rommem[19416] <= 16'hFFFF;
rommem[19417] <= 16'hFFFF;
rommem[19418] <= 16'hFFFF;
rommem[19419] <= 16'hFFFF;
rommem[19420] <= 16'hFFFF;
rommem[19421] <= 16'hFFFF;
rommem[19422] <= 16'hFFFF;
rommem[19423] <= 16'hFFFF;
rommem[19424] <= 16'hFFFF;
rommem[19425] <= 16'hFFFF;
rommem[19426] <= 16'hFFFF;
rommem[19427] <= 16'hFFFF;
rommem[19428] <= 16'hFFFF;
rommem[19429] <= 16'hFFFF;
rommem[19430] <= 16'hFFFF;
rommem[19431] <= 16'hFFFF;
rommem[19432] <= 16'hFFFF;
rommem[19433] <= 16'hFFFF;
rommem[19434] <= 16'hFFFF;
rommem[19435] <= 16'hFFFF;
rommem[19436] <= 16'hFFFF;
rommem[19437] <= 16'hFFFF;
rommem[19438] <= 16'hFFFF;
rommem[19439] <= 16'hFFFF;
rommem[19440] <= 16'hFFFF;
rommem[19441] <= 16'hFFFF;
rommem[19442] <= 16'hFFFF;
rommem[19443] <= 16'hFFFF;
rommem[19444] <= 16'hFFFF;
rommem[19445] <= 16'hFFFF;
rommem[19446] <= 16'hFFFF;
rommem[19447] <= 16'hFFFF;
rommem[19448] <= 16'hFFFF;
rommem[19449] <= 16'hFFFF;
rommem[19450] <= 16'hFFFF;
rommem[19451] <= 16'hFFFF;
rommem[19452] <= 16'hFFFF;
rommem[19453] <= 16'hFFFF;
rommem[19454] <= 16'hFFFF;
rommem[19455] <= 16'hFFFF;
rommem[19456] <= 16'hFFFF;
rommem[19457] <= 16'hFFFF;
rommem[19458] <= 16'hFFFF;
rommem[19459] <= 16'hFFFF;
rommem[19460] <= 16'hFFFF;
rommem[19461] <= 16'hFFFF;
rommem[19462] <= 16'hFFFF;
rommem[19463] <= 16'hFFFF;
rommem[19464] <= 16'hFFFF;
rommem[19465] <= 16'hFFFF;
rommem[19466] <= 16'hFFFF;
rommem[19467] <= 16'hFFFF;
rommem[19468] <= 16'hFFFF;
rommem[19469] <= 16'hFFFF;
rommem[19470] <= 16'hFFFF;
rommem[19471] <= 16'hFFFF;
rommem[19472] <= 16'hFFFF;
rommem[19473] <= 16'hFFFF;
rommem[19474] <= 16'hFFFF;
rommem[19475] <= 16'hFFFF;
rommem[19476] <= 16'hFFFF;
rommem[19477] <= 16'hFFFF;
rommem[19478] <= 16'hFFFF;
rommem[19479] <= 16'hFFFF;
rommem[19480] <= 16'hFFFF;
rommem[19481] <= 16'hFFFF;
rommem[19482] <= 16'hFFFF;
rommem[19483] <= 16'hFFFF;
rommem[19484] <= 16'hFFFF;
rommem[19485] <= 16'hFFFF;
rommem[19486] <= 16'hFFFF;
rommem[19487] <= 16'hFFFF;
rommem[19488] <= 16'hFFFF;
rommem[19489] <= 16'hFFFF;
rommem[19490] <= 16'hFFFF;
rommem[19491] <= 16'hFFFF;
rommem[19492] <= 16'hFFFF;
rommem[19493] <= 16'hFFFF;
rommem[19494] <= 16'hFFFF;
rommem[19495] <= 16'hFFFF;
rommem[19496] <= 16'hFFFF;
rommem[19497] <= 16'hFFFF;
rommem[19498] <= 16'hFFFF;
rommem[19499] <= 16'hFFFF;
rommem[19500] <= 16'hFFFF;
rommem[19501] <= 16'hFFFF;
rommem[19502] <= 16'hFFFF;
rommem[19503] <= 16'hFFFF;
rommem[19504] <= 16'hFFFF;
rommem[19505] <= 16'hFFFF;
rommem[19506] <= 16'hFFFF;
rommem[19507] <= 16'hFFFF;
rommem[19508] <= 16'hFFFF;
rommem[19509] <= 16'hFFFF;
rommem[19510] <= 16'hFFFF;
rommem[19511] <= 16'hFFFF;
rommem[19512] <= 16'hFFFF;
rommem[19513] <= 16'hFFFF;
rommem[19514] <= 16'hFFFF;
rommem[19515] <= 16'hFFFF;
rommem[19516] <= 16'hFFFF;
rommem[19517] <= 16'hFFFF;
rommem[19518] <= 16'hFFFF;
rommem[19519] <= 16'hFFFF;
rommem[19520] <= 16'hFFFF;
rommem[19521] <= 16'hFFFF;
rommem[19522] <= 16'hFFFF;
rommem[19523] <= 16'hFFFF;
rommem[19524] <= 16'hFFFF;
rommem[19525] <= 16'hFFFF;
rommem[19526] <= 16'hFFFF;
rommem[19527] <= 16'hFFFF;
rommem[19528] <= 16'hFFFF;
rommem[19529] <= 16'hFFFF;
rommem[19530] <= 16'hFFFF;
rommem[19531] <= 16'hFFFF;
rommem[19532] <= 16'hFFFF;
rommem[19533] <= 16'hFFFF;
rommem[19534] <= 16'hFFFF;
rommem[19535] <= 16'hFFFF;
rommem[19536] <= 16'hFFFF;
rommem[19537] <= 16'hFFFF;
rommem[19538] <= 16'hFFFF;
rommem[19539] <= 16'hFFFF;
rommem[19540] <= 16'hFFFF;
rommem[19541] <= 16'hFFFF;
rommem[19542] <= 16'hFFFF;
rommem[19543] <= 16'hFFFF;
rommem[19544] <= 16'hFFFF;
rommem[19545] <= 16'hFFFF;
rommem[19546] <= 16'hFFFF;
rommem[19547] <= 16'hFFFF;
rommem[19548] <= 16'hFFFF;
rommem[19549] <= 16'hFFFF;
rommem[19550] <= 16'hFFFF;
rommem[19551] <= 16'hFFFF;
rommem[19552] <= 16'hFFFF;
rommem[19553] <= 16'hFFFF;
rommem[19554] <= 16'hFFFF;
rommem[19555] <= 16'hFFFF;
rommem[19556] <= 16'hFFFF;
rommem[19557] <= 16'hFFFF;
rommem[19558] <= 16'hFFFF;
rommem[19559] <= 16'hFFFF;
rommem[19560] <= 16'hFFFF;
rommem[19561] <= 16'hFFFF;
rommem[19562] <= 16'hFFFF;
rommem[19563] <= 16'hFFFF;
rommem[19564] <= 16'hFFFF;
rommem[19565] <= 16'hFFFF;
rommem[19566] <= 16'hFFFF;
rommem[19567] <= 16'hFFFF;
rommem[19568] <= 16'hFFFF;
rommem[19569] <= 16'hFFFF;
rommem[19570] <= 16'hFFFF;
rommem[19571] <= 16'hFFFF;
rommem[19572] <= 16'hFFFF;
rommem[19573] <= 16'hFFFF;
rommem[19574] <= 16'hFFFF;
rommem[19575] <= 16'hFFFF;
rommem[19576] <= 16'hFFFF;
rommem[19577] <= 16'hFFFF;
rommem[19578] <= 16'hFFFF;
rommem[19579] <= 16'hFFFF;
rommem[19580] <= 16'hFFFF;
rommem[19581] <= 16'hFFFF;
rommem[19582] <= 16'hFFFF;
rommem[19583] <= 16'hFFFF;
rommem[19584] <= 16'hFFFF;
rommem[19585] <= 16'hFFFF;
rommem[19586] <= 16'hFFFF;
rommem[19587] <= 16'hFFFF;
rommem[19588] <= 16'hFFFF;
rommem[19589] <= 16'hFFFF;
rommem[19590] <= 16'hFFFF;
rommem[19591] <= 16'hFFFF;
rommem[19592] <= 16'hFFFF;
rommem[19593] <= 16'hFFFF;
rommem[19594] <= 16'hFFFF;
rommem[19595] <= 16'hFFFF;
rommem[19596] <= 16'hFFFF;
rommem[19597] <= 16'hFFFF;
rommem[19598] <= 16'hFFFF;
rommem[19599] <= 16'hFFFF;
rommem[19600] <= 16'hFFFF;
rommem[19601] <= 16'hFFFF;
rommem[19602] <= 16'hFFFF;
rommem[19603] <= 16'hFFFF;
rommem[19604] <= 16'hFFFF;
rommem[19605] <= 16'hFFFF;
rommem[19606] <= 16'hFFFF;
rommem[19607] <= 16'hFFFF;
rommem[19608] <= 16'hFFFF;
rommem[19609] <= 16'hFFFF;
rommem[19610] <= 16'hFFFF;
rommem[19611] <= 16'hFFFF;
rommem[19612] <= 16'hFFFF;
rommem[19613] <= 16'hFFFF;
rommem[19614] <= 16'hFFFF;
rommem[19615] <= 16'hFFFF;
rommem[19616] <= 16'hFFFF;
rommem[19617] <= 16'hFFFF;
rommem[19618] <= 16'hFFFF;
rommem[19619] <= 16'hFFFF;
rommem[19620] <= 16'hFFFF;
rommem[19621] <= 16'hFFFF;
rommem[19622] <= 16'hFFFF;
rommem[19623] <= 16'hFFFF;
rommem[19624] <= 16'hFFFF;
rommem[19625] <= 16'hFFFF;
rommem[19626] <= 16'hFFFF;
rommem[19627] <= 16'hFFFF;
rommem[19628] <= 16'hFFFF;
rommem[19629] <= 16'hFFFF;
rommem[19630] <= 16'hFFFF;
rommem[19631] <= 16'hFFFF;
rommem[19632] <= 16'hFFFF;
rommem[19633] <= 16'hFFFF;
rommem[19634] <= 16'hFFFF;
rommem[19635] <= 16'hFFFF;
rommem[19636] <= 16'hFFFF;
rommem[19637] <= 16'hFFFF;
rommem[19638] <= 16'hFFFF;
rommem[19639] <= 16'hFFFF;
rommem[19640] <= 16'hFFFF;
rommem[19641] <= 16'hFFFF;
rommem[19642] <= 16'hFFFF;
rommem[19643] <= 16'hFFFF;
rommem[19644] <= 16'hFFFF;
rommem[19645] <= 16'hFFFF;
rommem[19646] <= 16'hFFFF;
rommem[19647] <= 16'hFFFF;
rommem[19648] <= 16'hFFFF;
rommem[19649] <= 16'hFFFF;
rommem[19650] <= 16'hFFFF;
rommem[19651] <= 16'hFFFF;
rommem[19652] <= 16'hFFFF;
rommem[19653] <= 16'hFFFF;
rommem[19654] <= 16'hFFFF;
rommem[19655] <= 16'hFFFF;
rommem[19656] <= 16'hFFFF;
rommem[19657] <= 16'hFFFF;
rommem[19658] <= 16'hFFFF;
rommem[19659] <= 16'hFFFF;
rommem[19660] <= 16'hFFFF;
rommem[19661] <= 16'hFFFF;
rommem[19662] <= 16'hFFFF;
rommem[19663] <= 16'hFFFF;
rommem[19664] <= 16'hFFFF;
rommem[19665] <= 16'hFFFF;
rommem[19666] <= 16'hFFFF;
rommem[19667] <= 16'hFFFF;
rommem[19668] <= 16'hFFFF;
rommem[19669] <= 16'hFFFF;
rommem[19670] <= 16'hFFFF;
rommem[19671] <= 16'hFFFF;
rommem[19672] <= 16'hFFFF;
rommem[19673] <= 16'hFFFF;
rommem[19674] <= 16'hFFFF;
rommem[19675] <= 16'hFFFF;
rommem[19676] <= 16'hFFFF;
rommem[19677] <= 16'hFFFF;
rommem[19678] <= 16'hFFFF;
rommem[19679] <= 16'hFFFF;
rommem[19680] <= 16'hFFFF;
rommem[19681] <= 16'hFFFF;
rommem[19682] <= 16'hFFFF;
rommem[19683] <= 16'hFFFF;
rommem[19684] <= 16'hFFFF;
rommem[19685] <= 16'hFFFF;
rommem[19686] <= 16'hFFFF;
rommem[19687] <= 16'hFFFF;
rommem[19688] <= 16'hFFFF;
rommem[19689] <= 16'hFFFF;
rommem[19690] <= 16'hFFFF;
rommem[19691] <= 16'hFFFF;
rommem[19692] <= 16'hFFFF;
rommem[19693] <= 16'hFFFF;
rommem[19694] <= 16'hFFFF;
rommem[19695] <= 16'hFFFF;
rommem[19696] <= 16'hFFFF;
rommem[19697] <= 16'hFFFF;
rommem[19698] <= 16'hFFFF;
rommem[19699] <= 16'hFFFF;
rommem[19700] <= 16'hFFFF;
rommem[19701] <= 16'hFFFF;
rommem[19702] <= 16'hFFFF;
rommem[19703] <= 16'hFFFF;
rommem[19704] <= 16'hFFFF;
rommem[19705] <= 16'hFFFF;
rommem[19706] <= 16'hFFFF;
rommem[19707] <= 16'hFFFF;
rommem[19708] <= 16'hFFFF;
rommem[19709] <= 16'hFFFF;
rommem[19710] <= 16'hFFFF;
rommem[19711] <= 16'hFFFF;
rommem[19712] <= 16'hFFFF;
rommem[19713] <= 16'hFFFF;
rommem[19714] <= 16'hFFFF;
rommem[19715] <= 16'hFFFF;
rommem[19716] <= 16'hFFFF;
rommem[19717] <= 16'hFFFF;
rommem[19718] <= 16'hFFFF;
rommem[19719] <= 16'hFFFF;
rommem[19720] <= 16'hFFFF;
rommem[19721] <= 16'hFFFF;
rommem[19722] <= 16'hFFFF;
rommem[19723] <= 16'hFFFF;
rommem[19724] <= 16'hFFFF;
rommem[19725] <= 16'hFFFF;
rommem[19726] <= 16'hFFFF;
rommem[19727] <= 16'hFFFF;
rommem[19728] <= 16'hFFFF;
rommem[19729] <= 16'hFFFF;
rommem[19730] <= 16'hFFFF;
rommem[19731] <= 16'hFFFF;
rommem[19732] <= 16'hFFFF;
rommem[19733] <= 16'hFFFF;
rommem[19734] <= 16'hFFFF;
rommem[19735] <= 16'hFFFF;
rommem[19736] <= 16'hFFFF;
rommem[19737] <= 16'hFFFF;
rommem[19738] <= 16'hFFFF;
rommem[19739] <= 16'hFFFF;
rommem[19740] <= 16'hFFFF;
rommem[19741] <= 16'hFFFF;
rommem[19742] <= 16'hFFFF;
rommem[19743] <= 16'hFFFF;
rommem[19744] <= 16'hFFFF;
rommem[19745] <= 16'hFFFF;
rommem[19746] <= 16'hFFFF;
rommem[19747] <= 16'hFFFF;
rommem[19748] <= 16'hFFFF;
rommem[19749] <= 16'hFFFF;
rommem[19750] <= 16'hFFFF;
rommem[19751] <= 16'hFFFF;
rommem[19752] <= 16'hFFFF;
rommem[19753] <= 16'hFFFF;
rommem[19754] <= 16'hFFFF;
rommem[19755] <= 16'hFFFF;
rommem[19756] <= 16'hFFFF;
rommem[19757] <= 16'hFFFF;
rommem[19758] <= 16'hFFFF;
rommem[19759] <= 16'hFFFF;
rommem[19760] <= 16'hFFFF;
rommem[19761] <= 16'hFFFF;
rommem[19762] <= 16'hFFFF;
rommem[19763] <= 16'hFFFF;
rommem[19764] <= 16'hFFFF;
rommem[19765] <= 16'hFFFF;
rommem[19766] <= 16'hFFFF;
rommem[19767] <= 16'hFFFF;
rommem[19768] <= 16'hFFFF;
rommem[19769] <= 16'hFFFF;
rommem[19770] <= 16'hFFFF;
rommem[19771] <= 16'hFFFF;
rommem[19772] <= 16'hFFFF;
rommem[19773] <= 16'hFFFF;
rommem[19774] <= 16'hFFFF;
rommem[19775] <= 16'hFFFF;
rommem[19776] <= 16'hFFFF;
rommem[19777] <= 16'hFFFF;
rommem[19778] <= 16'hFFFF;
rommem[19779] <= 16'hFFFF;
rommem[19780] <= 16'hFFFF;
rommem[19781] <= 16'hFFFF;
rommem[19782] <= 16'hFFFF;
rommem[19783] <= 16'hFFFF;
rommem[19784] <= 16'hFFFF;
rommem[19785] <= 16'hFFFF;
rommem[19786] <= 16'hFFFF;
rommem[19787] <= 16'hFFFF;
rommem[19788] <= 16'hFFFF;
rommem[19789] <= 16'hFFFF;
rommem[19790] <= 16'hFFFF;
rommem[19791] <= 16'hFFFF;
rommem[19792] <= 16'hFFFF;
rommem[19793] <= 16'hFFFF;
rommem[19794] <= 16'hFFFF;
rommem[19795] <= 16'hFFFF;
rommem[19796] <= 16'hFFFF;
rommem[19797] <= 16'hFFFF;
rommem[19798] <= 16'hFFFF;
rommem[19799] <= 16'hFFFF;
rommem[19800] <= 16'hFFFF;
rommem[19801] <= 16'hFFFF;
rommem[19802] <= 16'hFFFF;
rommem[19803] <= 16'hFFFF;
rommem[19804] <= 16'hFFFF;
rommem[19805] <= 16'hFFFF;
rommem[19806] <= 16'hFFFF;
rommem[19807] <= 16'hFFFF;
rommem[19808] <= 16'hFFFF;
rommem[19809] <= 16'hFFFF;
rommem[19810] <= 16'hFFFF;
rommem[19811] <= 16'hFFFF;
rommem[19812] <= 16'hFFFF;
rommem[19813] <= 16'hFFFF;
rommem[19814] <= 16'hFFFF;
rommem[19815] <= 16'hFFFF;
rommem[19816] <= 16'hFFFF;
rommem[19817] <= 16'hFFFF;
rommem[19818] <= 16'hFFFF;
rommem[19819] <= 16'hFFFF;
rommem[19820] <= 16'hFFFF;
rommem[19821] <= 16'hFFFF;
rommem[19822] <= 16'hFFFF;
rommem[19823] <= 16'hFFFF;
rommem[19824] <= 16'hFFFF;
rommem[19825] <= 16'hFFFF;
rommem[19826] <= 16'hFFFF;
rommem[19827] <= 16'hFFFF;
rommem[19828] <= 16'hFFFF;
rommem[19829] <= 16'hFFFF;
rommem[19830] <= 16'hFFFF;
rommem[19831] <= 16'hFFFF;
rommem[19832] <= 16'hFFFF;
rommem[19833] <= 16'hFFFF;
rommem[19834] <= 16'hFFFF;
rommem[19835] <= 16'hFFFF;
rommem[19836] <= 16'hFFFF;
rommem[19837] <= 16'hFFFF;
rommem[19838] <= 16'hFFFF;
rommem[19839] <= 16'hFFFF;
rommem[19840] <= 16'hFFFF;
rommem[19841] <= 16'hFFFF;
rommem[19842] <= 16'hFFFF;
rommem[19843] <= 16'hFFFF;
rommem[19844] <= 16'hFFFF;
rommem[19845] <= 16'hFFFF;
rommem[19846] <= 16'hFFFF;
rommem[19847] <= 16'hFFFF;
rommem[19848] <= 16'hFFFF;
rommem[19849] <= 16'hFFFF;
rommem[19850] <= 16'hFFFF;
rommem[19851] <= 16'hFFFF;
rommem[19852] <= 16'hFFFF;
rommem[19853] <= 16'hFFFF;
rommem[19854] <= 16'hFFFF;
rommem[19855] <= 16'hFFFF;
rommem[19856] <= 16'hFFFF;
rommem[19857] <= 16'hFFFF;
rommem[19858] <= 16'hFFFF;
rommem[19859] <= 16'hFFFF;
rommem[19860] <= 16'hFFFF;
rommem[19861] <= 16'hFFFF;
rommem[19862] <= 16'hFFFF;
rommem[19863] <= 16'hFFFF;
rommem[19864] <= 16'hFFFF;
rommem[19865] <= 16'hFFFF;
rommem[19866] <= 16'hFFFF;
rommem[19867] <= 16'hFFFF;
rommem[19868] <= 16'hFFFF;
rommem[19869] <= 16'hFFFF;
rommem[19870] <= 16'hFFFF;
rommem[19871] <= 16'hFFFF;
rommem[19872] <= 16'hFFFF;
rommem[19873] <= 16'hFFFF;
rommem[19874] <= 16'hFFFF;
rommem[19875] <= 16'hFFFF;
rommem[19876] <= 16'hFFFF;
rommem[19877] <= 16'hFFFF;
rommem[19878] <= 16'hFFFF;
rommem[19879] <= 16'hFFFF;
rommem[19880] <= 16'hFFFF;
rommem[19881] <= 16'hFFFF;
rommem[19882] <= 16'hFFFF;
rommem[19883] <= 16'hFFFF;
rommem[19884] <= 16'hFFFF;
rommem[19885] <= 16'hFFFF;
rommem[19886] <= 16'hFFFF;
rommem[19887] <= 16'hFFFF;
rommem[19888] <= 16'hFFFF;
rommem[19889] <= 16'hFFFF;
rommem[19890] <= 16'hFFFF;
rommem[19891] <= 16'hFFFF;
rommem[19892] <= 16'hFFFF;
rommem[19893] <= 16'hFFFF;
rommem[19894] <= 16'hFFFF;
rommem[19895] <= 16'hFFFF;
rommem[19896] <= 16'hFFFF;
rommem[19897] <= 16'hFFFF;
rommem[19898] <= 16'hFFFF;
rommem[19899] <= 16'hFFFF;
rommem[19900] <= 16'hFFFF;
rommem[19901] <= 16'hFFFF;
rommem[19902] <= 16'hFFFF;
rommem[19903] <= 16'hFFFF;
rommem[19904] <= 16'hFFFF;
rommem[19905] <= 16'hFFFF;
rommem[19906] <= 16'hFFFF;
rommem[19907] <= 16'hFFFF;
rommem[19908] <= 16'hFFFF;
rommem[19909] <= 16'hFFFF;
rommem[19910] <= 16'hFFFF;
rommem[19911] <= 16'hFFFF;
rommem[19912] <= 16'hFFFF;
rommem[19913] <= 16'hFFFF;
rommem[19914] <= 16'hFFFF;
rommem[19915] <= 16'hFFFF;
rommem[19916] <= 16'hFFFF;
rommem[19917] <= 16'hFFFF;
rommem[19918] <= 16'hFFFF;
rommem[19919] <= 16'hFFFF;
rommem[19920] <= 16'hFFFF;
rommem[19921] <= 16'hFFFF;
rommem[19922] <= 16'hFFFF;
rommem[19923] <= 16'hFFFF;
rommem[19924] <= 16'hFFFF;
rommem[19925] <= 16'hFFFF;
rommem[19926] <= 16'hFFFF;
rommem[19927] <= 16'hFFFF;
rommem[19928] <= 16'hFFFF;
rommem[19929] <= 16'hFFFF;
rommem[19930] <= 16'hFFFF;
rommem[19931] <= 16'hFFFF;
rommem[19932] <= 16'hFFFF;
rommem[19933] <= 16'hFFFF;
rommem[19934] <= 16'hFFFF;
rommem[19935] <= 16'hFFFF;
rommem[19936] <= 16'hFFFF;
rommem[19937] <= 16'hFFFF;
rommem[19938] <= 16'hFFFF;
rommem[19939] <= 16'hFFFF;
rommem[19940] <= 16'hFFFF;
rommem[19941] <= 16'hFFFF;
rommem[19942] <= 16'hFFFF;
rommem[19943] <= 16'hFFFF;
rommem[19944] <= 16'hFFFF;
rommem[19945] <= 16'hFFFF;
rommem[19946] <= 16'hFFFF;
rommem[19947] <= 16'hFFFF;
rommem[19948] <= 16'hFFFF;
rommem[19949] <= 16'hFFFF;
rommem[19950] <= 16'hFFFF;
rommem[19951] <= 16'hFFFF;
rommem[19952] <= 16'hFFFF;
rommem[19953] <= 16'hFFFF;
rommem[19954] <= 16'hFFFF;
rommem[19955] <= 16'hFFFF;
rommem[19956] <= 16'hFFFF;
rommem[19957] <= 16'hFFFF;
rommem[19958] <= 16'hFFFF;
rommem[19959] <= 16'hFFFF;
rommem[19960] <= 16'hFFFF;
rommem[19961] <= 16'hFFFF;
rommem[19962] <= 16'hFFFF;
rommem[19963] <= 16'hFFFF;
rommem[19964] <= 16'hFFFF;
rommem[19965] <= 16'hFFFF;
rommem[19966] <= 16'hFFFF;
rommem[19967] <= 16'hFFFF;
rommem[19968] <= 16'hFFFF;
rommem[19969] <= 16'hFFFF;
rommem[19970] <= 16'hFFFF;
rommem[19971] <= 16'hFFFF;
rommem[19972] <= 16'hFFFF;
rommem[19973] <= 16'hFFFF;
rommem[19974] <= 16'hFFFF;
rommem[19975] <= 16'hFFFF;
rommem[19976] <= 16'hFFFF;
rommem[19977] <= 16'hFFFF;
rommem[19978] <= 16'hFFFF;
rommem[19979] <= 16'hFFFF;
rommem[19980] <= 16'hFFFF;
rommem[19981] <= 16'hFFFF;
rommem[19982] <= 16'hFFFF;
rommem[19983] <= 16'hFFFF;
rommem[19984] <= 16'hFFFF;
rommem[19985] <= 16'hFFFF;
rommem[19986] <= 16'hFFFF;
rommem[19987] <= 16'hFFFF;
rommem[19988] <= 16'hFFFF;
rommem[19989] <= 16'hFFFF;
rommem[19990] <= 16'hFFFF;
rommem[19991] <= 16'hFFFF;
rommem[19992] <= 16'hFFFF;
rommem[19993] <= 16'hFFFF;
rommem[19994] <= 16'hFFFF;
rommem[19995] <= 16'hFFFF;
rommem[19996] <= 16'hFFFF;
rommem[19997] <= 16'hFFFF;
rommem[19998] <= 16'hFFFF;
rommem[19999] <= 16'hFFFF;
rommem[20000] <= 16'hFFFF;
rommem[20001] <= 16'hFFFF;
rommem[20002] <= 16'hFFFF;
rommem[20003] <= 16'hFFFF;
rommem[20004] <= 16'hFFFF;
rommem[20005] <= 16'hFFFF;
rommem[20006] <= 16'hFFFF;
rommem[20007] <= 16'hFFFF;
rommem[20008] <= 16'hFFFF;
rommem[20009] <= 16'hFFFF;
rommem[20010] <= 16'hFFFF;
rommem[20011] <= 16'hFFFF;
rommem[20012] <= 16'hFFFF;
rommem[20013] <= 16'hFFFF;
rommem[20014] <= 16'hFFFF;
rommem[20015] <= 16'hFFFF;
rommem[20016] <= 16'hFFFF;
rommem[20017] <= 16'hFFFF;
rommem[20018] <= 16'hFFFF;
rommem[20019] <= 16'hFFFF;
rommem[20020] <= 16'hFFFF;
rommem[20021] <= 16'hFFFF;
rommem[20022] <= 16'hFFFF;
rommem[20023] <= 16'hFFFF;
rommem[20024] <= 16'hFFFF;
rommem[20025] <= 16'hFFFF;
rommem[20026] <= 16'hFFFF;
rommem[20027] <= 16'hFFFF;
rommem[20028] <= 16'hFFFF;
rommem[20029] <= 16'hFFFF;
rommem[20030] <= 16'hFFFF;
rommem[20031] <= 16'hFFFF;
rommem[20032] <= 16'hFFFF;
rommem[20033] <= 16'hFFFF;
rommem[20034] <= 16'hFFFF;
rommem[20035] <= 16'hFFFF;
rommem[20036] <= 16'hFFFF;
rommem[20037] <= 16'hFFFF;
rommem[20038] <= 16'hFFFF;
rommem[20039] <= 16'hFFFF;
rommem[20040] <= 16'hFFFF;
rommem[20041] <= 16'hFFFF;
rommem[20042] <= 16'hFFFF;
rommem[20043] <= 16'hFFFF;
rommem[20044] <= 16'hFFFF;
rommem[20045] <= 16'hFFFF;
rommem[20046] <= 16'hFFFF;
rommem[20047] <= 16'hFFFF;
rommem[20048] <= 16'hFFFF;
rommem[20049] <= 16'hFFFF;
rommem[20050] <= 16'hFFFF;
rommem[20051] <= 16'hFFFF;
rommem[20052] <= 16'hFFFF;
rommem[20053] <= 16'hFFFF;
rommem[20054] <= 16'hFFFF;
rommem[20055] <= 16'hFFFF;
rommem[20056] <= 16'hFFFF;
rommem[20057] <= 16'hFFFF;
rommem[20058] <= 16'hFFFF;
rommem[20059] <= 16'hFFFF;
rommem[20060] <= 16'hFFFF;
rommem[20061] <= 16'hFFFF;
rommem[20062] <= 16'hFFFF;
rommem[20063] <= 16'hFFFF;
rommem[20064] <= 16'hFFFF;
rommem[20065] <= 16'hFFFF;
rommem[20066] <= 16'hFFFF;
rommem[20067] <= 16'hFFFF;
rommem[20068] <= 16'hFFFF;
rommem[20069] <= 16'hFFFF;
rommem[20070] <= 16'hFFFF;
rommem[20071] <= 16'hFFFF;
rommem[20072] <= 16'hFFFF;
rommem[20073] <= 16'hFFFF;
rommem[20074] <= 16'hFFFF;
rommem[20075] <= 16'hFFFF;
rommem[20076] <= 16'hFFFF;
rommem[20077] <= 16'hFFFF;
rommem[20078] <= 16'hFFFF;
rommem[20079] <= 16'hFFFF;
rommem[20080] <= 16'hFFFF;
rommem[20081] <= 16'hFFFF;
rommem[20082] <= 16'hFFFF;
rommem[20083] <= 16'hFFFF;
rommem[20084] <= 16'hFFFF;
rommem[20085] <= 16'hFFFF;
rommem[20086] <= 16'hFFFF;
rommem[20087] <= 16'hFFFF;
rommem[20088] <= 16'hFFFF;
rommem[20089] <= 16'hFFFF;
rommem[20090] <= 16'hFFFF;
rommem[20091] <= 16'hFFFF;
rommem[20092] <= 16'hFFFF;
rommem[20093] <= 16'hFFFF;
rommem[20094] <= 16'hFFFF;
rommem[20095] <= 16'hFFFF;
rommem[20096] <= 16'hFFFF;
rommem[20097] <= 16'hFFFF;
rommem[20098] <= 16'hFFFF;
rommem[20099] <= 16'hFFFF;
rommem[20100] <= 16'hFFFF;
rommem[20101] <= 16'hFFFF;
rommem[20102] <= 16'hFFFF;
rommem[20103] <= 16'hFFFF;
rommem[20104] <= 16'hFFFF;
rommem[20105] <= 16'hFFFF;
rommem[20106] <= 16'hFFFF;
rommem[20107] <= 16'hFFFF;
rommem[20108] <= 16'hFFFF;
rommem[20109] <= 16'hFFFF;
rommem[20110] <= 16'hFFFF;
rommem[20111] <= 16'hFFFF;
rommem[20112] <= 16'hFFFF;
rommem[20113] <= 16'hFFFF;
rommem[20114] <= 16'hFFFF;
rommem[20115] <= 16'hFFFF;
rommem[20116] <= 16'hFFFF;
rommem[20117] <= 16'hFFFF;
rommem[20118] <= 16'hFFFF;
rommem[20119] <= 16'hFFFF;
rommem[20120] <= 16'hFFFF;
rommem[20121] <= 16'hFFFF;
rommem[20122] <= 16'hFFFF;
rommem[20123] <= 16'hFFFF;
rommem[20124] <= 16'hFFFF;
rommem[20125] <= 16'hFFFF;
rommem[20126] <= 16'hFFFF;
rommem[20127] <= 16'hFFFF;
rommem[20128] <= 16'hFFFF;
rommem[20129] <= 16'hFFFF;
rommem[20130] <= 16'hFFFF;
rommem[20131] <= 16'hFFFF;
rommem[20132] <= 16'hFFFF;
rommem[20133] <= 16'hFFFF;
rommem[20134] <= 16'hFFFF;
rommem[20135] <= 16'hFFFF;
rommem[20136] <= 16'hFFFF;
rommem[20137] <= 16'hFFFF;
rommem[20138] <= 16'hFFFF;
rommem[20139] <= 16'hFFFF;
rommem[20140] <= 16'hFFFF;
rommem[20141] <= 16'hFFFF;
rommem[20142] <= 16'hFFFF;
rommem[20143] <= 16'hFFFF;
rommem[20144] <= 16'hFFFF;
rommem[20145] <= 16'hFFFF;
rommem[20146] <= 16'hFFFF;
rommem[20147] <= 16'hFFFF;
rommem[20148] <= 16'hFFFF;
rommem[20149] <= 16'hFFFF;
rommem[20150] <= 16'hFFFF;
rommem[20151] <= 16'hFFFF;
rommem[20152] <= 16'hFFFF;
rommem[20153] <= 16'hFFFF;
rommem[20154] <= 16'hFFFF;
rommem[20155] <= 16'hFFFF;
rommem[20156] <= 16'hFFFF;
rommem[20157] <= 16'hFFFF;
rommem[20158] <= 16'hFFFF;
rommem[20159] <= 16'hFFFF;
rommem[20160] <= 16'hFFFF;
rommem[20161] <= 16'hFFFF;
rommem[20162] <= 16'hFFFF;
rommem[20163] <= 16'hFFFF;
rommem[20164] <= 16'hFFFF;
rommem[20165] <= 16'hFFFF;
rommem[20166] <= 16'hFFFF;
rommem[20167] <= 16'hFFFF;
rommem[20168] <= 16'hFFFF;
rommem[20169] <= 16'hFFFF;
rommem[20170] <= 16'hFFFF;
rommem[20171] <= 16'hFFFF;
rommem[20172] <= 16'hFFFF;
rommem[20173] <= 16'hFFFF;
rommem[20174] <= 16'hFFFF;
rommem[20175] <= 16'hFFFF;
rommem[20176] <= 16'hFFFF;
rommem[20177] <= 16'hFFFF;
rommem[20178] <= 16'hFFFF;
rommem[20179] <= 16'hFFFF;
rommem[20180] <= 16'hFFFF;
rommem[20181] <= 16'hFFFF;
rommem[20182] <= 16'hFFFF;
rommem[20183] <= 16'hFFFF;
rommem[20184] <= 16'hFFFF;
rommem[20185] <= 16'hFFFF;
rommem[20186] <= 16'hFFFF;
rommem[20187] <= 16'hFFFF;
rommem[20188] <= 16'hFFFF;
rommem[20189] <= 16'hFFFF;
rommem[20190] <= 16'hFFFF;
rommem[20191] <= 16'hFFFF;
rommem[20192] <= 16'hFFFF;
rommem[20193] <= 16'hFFFF;
rommem[20194] <= 16'hFFFF;
rommem[20195] <= 16'hFFFF;
rommem[20196] <= 16'hFFFF;
rommem[20197] <= 16'hFFFF;
rommem[20198] <= 16'hFFFF;
rommem[20199] <= 16'hFFFF;
rommem[20200] <= 16'hFFFF;
rommem[20201] <= 16'hFFFF;
rommem[20202] <= 16'hFFFF;
rommem[20203] <= 16'hFFFF;
rommem[20204] <= 16'hFFFF;
rommem[20205] <= 16'hFFFF;
rommem[20206] <= 16'hFFFF;
rommem[20207] <= 16'hFFFF;
rommem[20208] <= 16'hFFFF;
rommem[20209] <= 16'hFFFF;
rommem[20210] <= 16'hFFFF;
rommem[20211] <= 16'hFFFF;
rommem[20212] <= 16'hFFFF;
rommem[20213] <= 16'hFFFF;
rommem[20214] <= 16'hFFFF;
rommem[20215] <= 16'hFFFF;
rommem[20216] <= 16'hFFFF;
rommem[20217] <= 16'hFFFF;
rommem[20218] <= 16'hFFFF;
rommem[20219] <= 16'hFFFF;
rommem[20220] <= 16'hFFFF;
rommem[20221] <= 16'hFFFF;
rommem[20222] <= 16'hFFFF;
rommem[20223] <= 16'hFFFF;
rommem[20224] <= 16'hFFFF;
rommem[20225] <= 16'hFFFF;
rommem[20226] <= 16'hFFFF;
rommem[20227] <= 16'hFFFF;
rommem[20228] <= 16'hFFFF;
rommem[20229] <= 16'hFFFF;
rommem[20230] <= 16'hFFFF;
rommem[20231] <= 16'hFFFF;
rommem[20232] <= 16'hFFFF;
rommem[20233] <= 16'hFFFF;
rommem[20234] <= 16'hFFFF;
rommem[20235] <= 16'hFFFF;
rommem[20236] <= 16'hFFFF;
rommem[20237] <= 16'hFFFF;
rommem[20238] <= 16'hFFFF;
rommem[20239] <= 16'hFFFF;
rommem[20240] <= 16'hFFFF;
rommem[20241] <= 16'hFFFF;
rommem[20242] <= 16'hFFFF;
rommem[20243] <= 16'hFFFF;
rommem[20244] <= 16'hFFFF;
rommem[20245] <= 16'hFFFF;
rommem[20246] <= 16'hFFFF;
rommem[20247] <= 16'hFFFF;
rommem[20248] <= 16'hFFFF;
rommem[20249] <= 16'hFFFF;
rommem[20250] <= 16'hFFFF;
rommem[20251] <= 16'hFFFF;
rommem[20252] <= 16'hFFFF;
rommem[20253] <= 16'hFFFF;
rommem[20254] <= 16'hFFFF;
rommem[20255] <= 16'hFFFF;
rommem[20256] <= 16'hFFFF;
rommem[20257] <= 16'hFFFF;
rommem[20258] <= 16'hFFFF;
rommem[20259] <= 16'hFFFF;
rommem[20260] <= 16'hFFFF;
rommem[20261] <= 16'hFFFF;
rommem[20262] <= 16'hFFFF;
rommem[20263] <= 16'hFFFF;
rommem[20264] <= 16'hFFFF;
rommem[20265] <= 16'hFFFF;
rommem[20266] <= 16'hFFFF;
rommem[20267] <= 16'hFFFF;
rommem[20268] <= 16'hFFFF;
rommem[20269] <= 16'hFFFF;
rommem[20270] <= 16'hFFFF;
rommem[20271] <= 16'hFFFF;
rommem[20272] <= 16'hFFFF;
rommem[20273] <= 16'hFFFF;
rommem[20274] <= 16'hFFFF;
rommem[20275] <= 16'hFFFF;
rommem[20276] <= 16'hFFFF;
rommem[20277] <= 16'hFFFF;
rommem[20278] <= 16'hFFFF;
rommem[20279] <= 16'hFFFF;
rommem[20280] <= 16'hFFFF;
rommem[20281] <= 16'hFFFF;
rommem[20282] <= 16'hFFFF;
rommem[20283] <= 16'hFFFF;
rommem[20284] <= 16'hFFFF;
rommem[20285] <= 16'hFFFF;
rommem[20286] <= 16'hFFFF;
rommem[20287] <= 16'hFFFF;
rommem[20288] <= 16'hFFFF;
rommem[20289] <= 16'hFFFF;
rommem[20290] <= 16'hFFFF;
rommem[20291] <= 16'hFFFF;
rommem[20292] <= 16'hFFFF;
rommem[20293] <= 16'hFFFF;
rommem[20294] <= 16'hFFFF;
rommem[20295] <= 16'hFFFF;
rommem[20296] <= 16'hFFFF;
rommem[20297] <= 16'hFFFF;
rommem[20298] <= 16'hFFFF;
rommem[20299] <= 16'hFFFF;
rommem[20300] <= 16'hFFFF;
rommem[20301] <= 16'hFFFF;
rommem[20302] <= 16'hFFFF;
rommem[20303] <= 16'hFFFF;
rommem[20304] <= 16'hFFFF;
rommem[20305] <= 16'hFFFF;
rommem[20306] <= 16'hFFFF;
rommem[20307] <= 16'hFFFF;
rommem[20308] <= 16'hFFFF;
rommem[20309] <= 16'hFFFF;
rommem[20310] <= 16'hFFFF;
rommem[20311] <= 16'hFFFF;
rommem[20312] <= 16'hFFFF;
rommem[20313] <= 16'hFFFF;
rommem[20314] <= 16'hFFFF;
rommem[20315] <= 16'hFFFF;
rommem[20316] <= 16'hFFFF;
rommem[20317] <= 16'hFFFF;
rommem[20318] <= 16'hFFFF;
rommem[20319] <= 16'hFFFF;
rommem[20320] <= 16'hFFFF;
rommem[20321] <= 16'hFFFF;
rommem[20322] <= 16'hFFFF;
rommem[20323] <= 16'hFFFF;
rommem[20324] <= 16'hFFFF;
rommem[20325] <= 16'hFFFF;
rommem[20326] <= 16'hFFFF;
rommem[20327] <= 16'hFFFF;
rommem[20328] <= 16'hFFFF;
rommem[20329] <= 16'hFFFF;
rommem[20330] <= 16'hFFFF;
rommem[20331] <= 16'hFFFF;
rommem[20332] <= 16'hFFFF;
rommem[20333] <= 16'hFFFF;
rommem[20334] <= 16'hFFFF;
rommem[20335] <= 16'hFFFF;
rommem[20336] <= 16'hFFFF;
rommem[20337] <= 16'hFFFF;
rommem[20338] <= 16'hFFFF;
rommem[20339] <= 16'hFFFF;
rommem[20340] <= 16'hFFFF;
rommem[20341] <= 16'hFFFF;
rommem[20342] <= 16'hFFFF;
rommem[20343] <= 16'hFFFF;
rommem[20344] <= 16'hFFFF;
rommem[20345] <= 16'hFFFF;
rommem[20346] <= 16'hFFFF;
rommem[20347] <= 16'hFFFF;
rommem[20348] <= 16'hFFFF;
rommem[20349] <= 16'hFFFF;
rommem[20350] <= 16'hFFFF;
rommem[20351] <= 16'hFFFF;
rommem[20352] <= 16'hFFFF;
rommem[20353] <= 16'hFFFF;
rommem[20354] <= 16'hFFFF;
rommem[20355] <= 16'hFFFF;
rommem[20356] <= 16'hFFFF;
rommem[20357] <= 16'hFFFF;
rommem[20358] <= 16'hFFFF;
rommem[20359] <= 16'hFFFF;
rommem[20360] <= 16'hFFFF;
rommem[20361] <= 16'hFFFF;
rommem[20362] <= 16'hFFFF;
rommem[20363] <= 16'hFFFF;
rommem[20364] <= 16'hFFFF;
rommem[20365] <= 16'hFFFF;
rommem[20366] <= 16'hFFFF;
rommem[20367] <= 16'hFFFF;
rommem[20368] <= 16'hFFFF;
rommem[20369] <= 16'hFFFF;
rommem[20370] <= 16'hFFFF;
rommem[20371] <= 16'hFFFF;
rommem[20372] <= 16'hFFFF;
rommem[20373] <= 16'hFFFF;
rommem[20374] <= 16'hFFFF;
rommem[20375] <= 16'hFFFF;
rommem[20376] <= 16'hFFFF;
rommem[20377] <= 16'hFFFF;
rommem[20378] <= 16'hFFFF;
rommem[20379] <= 16'hFFFF;
rommem[20380] <= 16'hFFFF;
rommem[20381] <= 16'hFFFF;
rommem[20382] <= 16'hFFFF;
rommem[20383] <= 16'hFFFF;
rommem[20384] <= 16'hFFFF;
rommem[20385] <= 16'hFFFF;
rommem[20386] <= 16'hFFFF;
rommem[20387] <= 16'hFFFF;
rommem[20388] <= 16'hFFFF;
rommem[20389] <= 16'hFFFF;
rommem[20390] <= 16'hFFFF;
rommem[20391] <= 16'hFFFF;
rommem[20392] <= 16'hFFFF;
rommem[20393] <= 16'hFFFF;
rommem[20394] <= 16'hFFFF;
rommem[20395] <= 16'hFFFF;
rommem[20396] <= 16'hFFFF;
rommem[20397] <= 16'hFFFF;
rommem[20398] <= 16'hFFFF;
rommem[20399] <= 16'hFFFF;
rommem[20400] <= 16'hFFFF;
rommem[20401] <= 16'hFFFF;
rommem[20402] <= 16'hFFFF;
rommem[20403] <= 16'hFFFF;
rommem[20404] <= 16'hFFFF;
rommem[20405] <= 16'hFFFF;
rommem[20406] <= 16'hFFFF;
rommem[20407] <= 16'hFFFF;
rommem[20408] <= 16'hFFFF;
rommem[20409] <= 16'hFFFF;
rommem[20410] <= 16'hFFFF;
rommem[20411] <= 16'hFFFF;
rommem[20412] <= 16'hFFFF;
rommem[20413] <= 16'hFFFF;
rommem[20414] <= 16'hFFFF;
rommem[20415] <= 16'hFFFF;
rommem[20416] <= 16'hFFFF;
rommem[20417] <= 16'hFFFF;
rommem[20418] <= 16'hFFFF;
rommem[20419] <= 16'hFFFF;
rommem[20420] <= 16'hFFFF;
rommem[20421] <= 16'hFFFF;
rommem[20422] <= 16'hFFFF;
rommem[20423] <= 16'hFFFF;
rommem[20424] <= 16'hFFFF;
rommem[20425] <= 16'hFFFF;
rommem[20426] <= 16'hFFFF;
rommem[20427] <= 16'hFFFF;
rommem[20428] <= 16'hFFFF;
rommem[20429] <= 16'hFFFF;
rommem[20430] <= 16'hFFFF;
rommem[20431] <= 16'hFFFF;
rommem[20432] <= 16'hFFFF;
rommem[20433] <= 16'hFFFF;
rommem[20434] <= 16'hFFFF;
rommem[20435] <= 16'hFFFF;
rommem[20436] <= 16'hFFFF;
rommem[20437] <= 16'hFFFF;
rommem[20438] <= 16'hFFFF;
rommem[20439] <= 16'hFFFF;
rommem[20440] <= 16'hFFFF;
rommem[20441] <= 16'hFFFF;
rommem[20442] <= 16'hFFFF;
rommem[20443] <= 16'hFFFF;
rommem[20444] <= 16'hFFFF;
rommem[20445] <= 16'hFFFF;
rommem[20446] <= 16'hFFFF;
rommem[20447] <= 16'hFFFF;
rommem[20448] <= 16'hFFFF;
rommem[20449] <= 16'hFFFF;
rommem[20450] <= 16'hFFFF;
rommem[20451] <= 16'hFFFF;
rommem[20452] <= 16'hFFFF;
rommem[20453] <= 16'hFFFF;
rommem[20454] <= 16'hFFFF;
rommem[20455] <= 16'hFFFF;
rommem[20456] <= 16'hFFFF;
rommem[20457] <= 16'hFFFF;
rommem[20458] <= 16'hFFFF;
rommem[20459] <= 16'hFFFF;
rommem[20460] <= 16'hFFFF;
rommem[20461] <= 16'hFFFF;
rommem[20462] <= 16'hFFFF;
rommem[20463] <= 16'hFFFF;
rommem[20464] <= 16'hFFFF;
rommem[20465] <= 16'hFFFF;
rommem[20466] <= 16'hFFFF;
rommem[20467] <= 16'hFFFF;
rommem[20468] <= 16'hFFFF;
rommem[20469] <= 16'hFFFF;
rommem[20470] <= 16'hFFFF;
rommem[20471] <= 16'hFFFF;
rommem[20472] <= 16'hFFFF;
rommem[20473] <= 16'hFFFF;
rommem[20474] <= 16'hFFFF;
rommem[20475] <= 16'hFFFF;
rommem[20476] <= 16'hFFFF;
rommem[20477] <= 16'hFFFF;
rommem[20478] <= 16'hFFFF;
rommem[20479] <= 16'hFFFF;
rommem[20480] <= 16'hFFFF;
rommem[20481] <= 16'hFFFF;
rommem[20482] <= 16'hFFFF;
rommem[20483] <= 16'hFFFF;
rommem[20484] <= 16'hFFFF;
rommem[20485] <= 16'hFFFF;
rommem[20486] <= 16'hFFFF;
rommem[20487] <= 16'hFFFF;
rommem[20488] <= 16'hFFFF;
rommem[20489] <= 16'hFFFF;
rommem[20490] <= 16'hFFFF;
rommem[20491] <= 16'hFFFF;
rommem[20492] <= 16'hFFFF;
rommem[20493] <= 16'hFFFF;
rommem[20494] <= 16'hFFFF;
rommem[20495] <= 16'hFFFF;
rommem[20496] <= 16'hFFFF;
rommem[20497] <= 16'hFFFF;
rommem[20498] <= 16'hFFFF;
rommem[20499] <= 16'hFFFF;
rommem[20500] <= 16'hFFFF;
rommem[20501] <= 16'hFFFF;
rommem[20502] <= 16'hFFFF;
rommem[20503] <= 16'hFFFF;
rommem[20504] <= 16'hFFFF;
rommem[20505] <= 16'hFFFF;
rommem[20506] <= 16'hFFFF;
rommem[20507] <= 16'hFFFF;
rommem[20508] <= 16'hFFFF;
rommem[20509] <= 16'hFFFF;
rommem[20510] <= 16'hFFFF;
rommem[20511] <= 16'hFFFF;
rommem[20512] <= 16'hFFFF;
rommem[20513] <= 16'hFFFF;
rommem[20514] <= 16'hFFFF;
rommem[20515] <= 16'hFFFF;
rommem[20516] <= 16'hFFFF;
rommem[20517] <= 16'hFFFF;
rommem[20518] <= 16'hFFFF;
rommem[20519] <= 16'hFFFF;
rommem[20520] <= 16'hFFFF;
rommem[20521] <= 16'hFFFF;
rommem[20522] <= 16'hFFFF;
rommem[20523] <= 16'hFFFF;
rommem[20524] <= 16'hFFFF;
rommem[20525] <= 16'hFFFF;
rommem[20526] <= 16'hFFFF;
rommem[20527] <= 16'hFFFF;
rommem[20528] <= 16'hFFFF;
rommem[20529] <= 16'hFFFF;
rommem[20530] <= 16'hFFFF;
rommem[20531] <= 16'hFFFF;
rommem[20532] <= 16'hFFFF;
rommem[20533] <= 16'hFFFF;
rommem[20534] <= 16'hFFFF;
rommem[20535] <= 16'hFFFF;
rommem[20536] <= 16'hFFFF;
rommem[20537] <= 16'hFFFF;
rommem[20538] <= 16'hFFFF;
rommem[20539] <= 16'hFFFF;
rommem[20540] <= 16'hFFFF;
rommem[20541] <= 16'hFFFF;
rommem[20542] <= 16'hFFFF;
rommem[20543] <= 16'hFFFF;
rommem[20544] <= 16'hFFFF;
rommem[20545] <= 16'hFFFF;
rommem[20546] <= 16'hFFFF;
rommem[20547] <= 16'hFFFF;
rommem[20548] <= 16'hFFFF;
rommem[20549] <= 16'hFFFF;
rommem[20550] <= 16'hFFFF;
rommem[20551] <= 16'hFFFF;
rommem[20552] <= 16'hFFFF;
rommem[20553] <= 16'hFFFF;
rommem[20554] <= 16'hFFFF;
rommem[20555] <= 16'hFFFF;
rommem[20556] <= 16'hFFFF;
rommem[20557] <= 16'hFFFF;
rommem[20558] <= 16'hFFFF;
rommem[20559] <= 16'hFFFF;
rommem[20560] <= 16'hFFFF;
rommem[20561] <= 16'hFFFF;
rommem[20562] <= 16'hFFFF;
rommem[20563] <= 16'hFFFF;
rommem[20564] <= 16'hFFFF;
rommem[20565] <= 16'hFFFF;
rommem[20566] <= 16'hFFFF;
rommem[20567] <= 16'hFFFF;
rommem[20568] <= 16'hFFFF;
rommem[20569] <= 16'hFFFF;
rommem[20570] <= 16'hFFFF;
rommem[20571] <= 16'hFFFF;
rommem[20572] <= 16'hFFFF;
rommem[20573] <= 16'hFFFF;
rommem[20574] <= 16'hFFFF;
rommem[20575] <= 16'hFFFF;
rommem[20576] <= 16'hFFFF;
rommem[20577] <= 16'hFFFF;
rommem[20578] <= 16'hFFFF;
rommem[20579] <= 16'hFFFF;
rommem[20580] <= 16'hFFFF;
rommem[20581] <= 16'hFFFF;
rommem[20582] <= 16'hFFFF;
rommem[20583] <= 16'hFFFF;
rommem[20584] <= 16'hFFFF;
rommem[20585] <= 16'hFFFF;
rommem[20586] <= 16'hFFFF;
rommem[20587] <= 16'hFFFF;
rommem[20588] <= 16'hFFFF;
rommem[20589] <= 16'hFFFF;
rommem[20590] <= 16'hFFFF;
rommem[20591] <= 16'hFFFF;
rommem[20592] <= 16'hFFFF;
rommem[20593] <= 16'hFFFF;
rommem[20594] <= 16'hFFFF;
rommem[20595] <= 16'hFFFF;
rommem[20596] <= 16'hFFFF;
rommem[20597] <= 16'hFFFF;
rommem[20598] <= 16'hFFFF;
rommem[20599] <= 16'hFFFF;
rommem[20600] <= 16'hFFFF;
rommem[20601] <= 16'hFFFF;
rommem[20602] <= 16'hFFFF;
rommem[20603] <= 16'hFFFF;
rommem[20604] <= 16'hFFFF;
rommem[20605] <= 16'hFFFF;
rommem[20606] <= 16'hFFFF;
rommem[20607] <= 16'hFFFF;
rommem[20608] <= 16'hFFFF;
rommem[20609] <= 16'hFFFF;
rommem[20610] <= 16'hFFFF;
rommem[20611] <= 16'hFFFF;
rommem[20612] <= 16'hFFFF;
rommem[20613] <= 16'hFFFF;
rommem[20614] <= 16'hFFFF;
rommem[20615] <= 16'hFFFF;
rommem[20616] <= 16'hFFFF;
rommem[20617] <= 16'hFFFF;
rommem[20618] <= 16'hFFFF;
rommem[20619] <= 16'hFFFF;
rommem[20620] <= 16'hFFFF;
rommem[20621] <= 16'hFFFF;
rommem[20622] <= 16'hFFFF;
rommem[20623] <= 16'hFFFF;
rommem[20624] <= 16'hFFFF;
rommem[20625] <= 16'hFFFF;
rommem[20626] <= 16'hFFFF;
rommem[20627] <= 16'hFFFF;
rommem[20628] <= 16'hFFFF;
rommem[20629] <= 16'hFFFF;
rommem[20630] <= 16'hFFFF;
rommem[20631] <= 16'hFFFF;
rommem[20632] <= 16'hFFFF;
rommem[20633] <= 16'hFFFF;
rommem[20634] <= 16'hFFFF;
rommem[20635] <= 16'hFFFF;
rommem[20636] <= 16'hFFFF;
rommem[20637] <= 16'hFFFF;
rommem[20638] <= 16'hFFFF;
rommem[20639] <= 16'hFFFF;
rommem[20640] <= 16'hFFFF;
rommem[20641] <= 16'hFFFF;
rommem[20642] <= 16'hFFFF;
rommem[20643] <= 16'hFFFF;
rommem[20644] <= 16'hFFFF;
rommem[20645] <= 16'hFFFF;
rommem[20646] <= 16'hFFFF;
rommem[20647] <= 16'hFFFF;
rommem[20648] <= 16'hFFFF;
rommem[20649] <= 16'hFFFF;
rommem[20650] <= 16'hFFFF;
rommem[20651] <= 16'hFFFF;
rommem[20652] <= 16'hFFFF;
rommem[20653] <= 16'hFFFF;
rommem[20654] <= 16'hFFFF;
rommem[20655] <= 16'hFFFF;
rommem[20656] <= 16'hFFFF;
rommem[20657] <= 16'hFFFF;
rommem[20658] <= 16'hFFFF;
rommem[20659] <= 16'hFFFF;
rommem[20660] <= 16'hFFFF;
rommem[20661] <= 16'hFFFF;
rommem[20662] <= 16'hFFFF;
rommem[20663] <= 16'hFFFF;
rommem[20664] <= 16'hFFFF;
rommem[20665] <= 16'hFFFF;
rommem[20666] <= 16'hFFFF;
rommem[20667] <= 16'hFFFF;
rommem[20668] <= 16'hFFFF;
rommem[20669] <= 16'hFFFF;
rommem[20670] <= 16'hFFFF;
rommem[20671] <= 16'hFFFF;
rommem[20672] <= 16'hFFFF;
rommem[20673] <= 16'hFFFF;
rommem[20674] <= 16'hFFFF;
rommem[20675] <= 16'hFFFF;
rommem[20676] <= 16'hFFFF;
rommem[20677] <= 16'hFFFF;
rommem[20678] <= 16'hFFFF;
rommem[20679] <= 16'hFFFF;
rommem[20680] <= 16'hFFFF;
rommem[20681] <= 16'hFFFF;
rommem[20682] <= 16'hFFFF;
rommem[20683] <= 16'hFFFF;
rommem[20684] <= 16'hFFFF;
rommem[20685] <= 16'hFFFF;
rommem[20686] <= 16'hFFFF;
rommem[20687] <= 16'hFFFF;
rommem[20688] <= 16'hFFFF;
rommem[20689] <= 16'hFFFF;
rommem[20690] <= 16'hFFFF;
rommem[20691] <= 16'hFFFF;
rommem[20692] <= 16'hFFFF;
rommem[20693] <= 16'hFFFF;
rommem[20694] <= 16'hFFFF;
rommem[20695] <= 16'hFFFF;
rommem[20696] <= 16'hFFFF;
rommem[20697] <= 16'hFFFF;
rommem[20698] <= 16'hFFFF;
rommem[20699] <= 16'hFFFF;
rommem[20700] <= 16'hFFFF;
rommem[20701] <= 16'hFFFF;
rommem[20702] <= 16'hFFFF;
rommem[20703] <= 16'hFFFF;
rommem[20704] <= 16'hFFFF;
rommem[20705] <= 16'hFFFF;
rommem[20706] <= 16'hFFFF;
rommem[20707] <= 16'hFFFF;
rommem[20708] <= 16'hFFFF;
rommem[20709] <= 16'hFFFF;
rommem[20710] <= 16'hFFFF;
rommem[20711] <= 16'hFFFF;
rommem[20712] <= 16'hFFFF;
rommem[20713] <= 16'hFFFF;
rommem[20714] <= 16'hFFFF;
rommem[20715] <= 16'hFFFF;
rommem[20716] <= 16'hFFFF;
rommem[20717] <= 16'hFFFF;
rommem[20718] <= 16'hFFFF;
rommem[20719] <= 16'hFFFF;
rommem[20720] <= 16'hFFFF;
rommem[20721] <= 16'hFFFF;
rommem[20722] <= 16'hFFFF;
rommem[20723] <= 16'hFFFF;
rommem[20724] <= 16'hFFFF;
rommem[20725] <= 16'hFFFF;
rommem[20726] <= 16'hFFFF;
rommem[20727] <= 16'hFFFF;
rommem[20728] <= 16'hFFFF;
rommem[20729] <= 16'hFFFF;
rommem[20730] <= 16'hFFFF;
rommem[20731] <= 16'hFFFF;
rommem[20732] <= 16'hFFFF;
rommem[20733] <= 16'hFFFF;
rommem[20734] <= 16'hFFFF;
rommem[20735] <= 16'hFFFF;
rommem[20736] <= 16'hFFFF;
rommem[20737] <= 16'hFFFF;
rommem[20738] <= 16'hFFFF;
rommem[20739] <= 16'hFFFF;
rommem[20740] <= 16'hFFFF;
rommem[20741] <= 16'hFFFF;
rommem[20742] <= 16'hFFFF;
rommem[20743] <= 16'hFFFF;
rommem[20744] <= 16'hFFFF;
rommem[20745] <= 16'hFFFF;
rommem[20746] <= 16'hFFFF;
rommem[20747] <= 16'hFFFF;
rommem[20748] <= 16'hFFFF;
rommem[20749] <= 16'hFFFF;
rommem[20750] <= 16'hFFFF;
rommem[20751] <= 16'hFFFF;
rommem[20752] <= 16'hFFFF;
rommem[20753] <= 16'hFFFF;
rommem[20754] <= 16'hFFFF;
rommem[20755] <= 16'hFFFF;
rommem[20756] <= 16'hFFFF;
rommem[20757] <= 16'hFFFF;
rommem[20758] <= 16'hFFFF;
rommem[20759] <= 16'hFFFF;
rommem[20760] <= 16'hFFFF;
rommem[20761] <= 16'hFFFF;
rommem[20762] <= 16'hFFFF;
rommem[20763] <= 16'hFFFF;
rommem[20764] <= 16'hFFFF;
rommem[20765] <= 16'hFFFF;
rommem[20766] <= 16'hFFFF;
rommem[20767] <= 16'hFFFF;
rommem[20768] <= 16'hFFFF;
rommem[20769] <= 16'hFFFF;
rommem[20770] <= 16'hFFFF;
rommem[20771] <= 16'hFFFF;
rommem[20772] <= 16'hFFFF;
rommem[20773] <= 16'hFFFF;
rommem[20774] <= 16'hFFFF;
rommem[20775] <= 16'hFFFF;
rommem[20776] <= 16'hFFFF;
rommem[20777] <= 16'hFFFF;
rommem[20778] <= 16'hFFFF;
rommem[20779] <= 16'hFFFF;
rommem[20780] <= 16'hFFFF;
rommem[20781] <= 16'hFFFF;
rommem[20782] <= 16'hFFFF;
rommem[20783] <= 16'hFFFF;
rommem[20784] <= 16'hFFFF;
rommem[20785] <= 16'hFFFF;
rommem[20786] <= 16'hFFFF;
rommem[20787] <= 16'hFFFF;
rommem[20788] <= 16'hFFFF;
rommem[20789] <= 16'hFFFF;
rommem[20790] <= 16'hFFFF;
rommem[20791] <= 16'hFFFF;
rommem[20792] <= 16'hFFFF;
rommem[20793] <= 16'hFFFF;
rommem[20794] <= 16'hFFFF;
rommem[20795] <= 16'hFFFF;
rommem[20796] <= 16'hFFFF;
rommem[20797] <= 16'hFFFF;
rommem[20798] <= 16'hFFFF;
rommem[20799] <= 16'hFFFF;
rommem[20800] <= 16'hFFFF;
rommem[20801] <= 16'hFFFF;
rommem[20802] <= 16'hFFFF;
rommem[20803] <= 16'hFFFF;
rommem[20804] <= 16'hFFFF;
rommem[20805] <= 16'hFFFF;
rommem[20806] <= 16'hFFFF;
rommem[20807] <= 16'hFFFF;
rommem[20808] <= 16'hFFFF;
rommem[20809] <= 16'hFFFF;
rommem[20810] <= 16'hFFFF;
rommem[20811] <= 16'hFFFF;
rommem[20812] <= 16'hFFFF;
rommem[20813] <= 16'hFFFF;
rommem[20814] <= 16'hFFFF;
rommem[20815] <= 16'hFFFF;
rommem[20816] <= 16'hFFFF;
rommem[20817] <= 16'hFFFF;
rommem[20818] <= 16'hFFFF;
rommem[20819] <= 16'hFFFF;
rommem[20820] <= 16'hFFFF;
rommem[20821] <= 16'hFFFF;
rommem[20822] <= 16'hFFFF;
rommem[20823] <= 16'hFFFF;
rommem[20824] <= 16'hFFFF;
rommem[20825] <= 16'hFFFF;
rommem[20826] <= 16'hFFFF;
rommem[20827] <= 16'hFFFF;
rommem[20828] <= 16'hFFFF;
rommem[20829] <= 16'hFFFF;
rommem[20830] <= 16'hFFFF;
rommem[20831] <= 16'hFFFF;
rommem[20832] <= 16'hFFFF;
rommem[20833] <= 16'hFFFF;
rommem[20834] <= 16'hFFFF;
rommem[20835] <= 16'hFFFF;
rommem[20836] <= 16'hFFFF;
rommem[20837] <= 16'hFFFF;
rommem[20838] <= 16'hFFFF;
rommem[20839] <= 16'hFFFF;
rommem[20840] <= 16'hFFFF;
rommem[20841] <= 16'hFFFF;
rommem[20842] <= 16'hFFFF;
rommem[20843] <= 16'hFFFF;
rommem[20844] <= 16'hFFFF;
rommem[20845] <= 16'hFFFF;
rommem[20846] <= 16'hFFFF;
rommem[20847] <= 16'hFFFF;
rommem[20848] <= 16'hFFFF;
rommem[20849] <= 16'hFFFF;
rommem[20850] <= 16'hFFFF;
rommem[20851] <= 16'hFFFF;
rommem[20852] <= 16'hFFFF;
rommem[20853] <= 16'hFFFF;
rommem[20854] <= 16'hFFFF;
rommem[20855] <= 16'hFFFF;
rommem[20856] <= 16'hFFFF;
rommem[20857] <= 16'hFFFF;
rommem[20858] <= 16'hFFFF;
rommem[20859] <= 16'hFFFF;
rommem[20860] <= 16'hFFFF;
rommem[20861] <= 16'hFFFF;
rommem[20862] <= 16'hFFFF;
rommem[20863] <= 16'hFFFF;
rommem[20864] <= 16'hFFFF;
rommem[20865] <= 16'hFFFF;
rommem[20866] <= 16'hFFFF;
rommem[20867] <= 16'hFFFF;
rommem[20868] <= 16'hFFFF;
rommem[20869] <= 16'hFFFF;
rommem[20870] <= 16'hFFFF;
rommem[20871] <= 16'hFFFF;
rommem[20872] <= 16'hFFFF;
rommem[20873] <= 16'hFFFF;
rommem[20874] <= 16'hFFFF;
rommem[20875] <= 16'hFFFF;
rommem[20876] <= 16'hFFFF;
rommem[20877] <= 16'hFFFF;
rommem[20878] <= 16'hFFFF;
rommem[20879] <= 16'hFFFF;
rommem[20880] <= 16'hFFFF;
rommem[20881] <= 16'hFFFF;
rommem[20882] <= 16'hFFFF;
rommem[20883] <= 16'hFFFF;
rommem[20884] <= 16'hFFFF;
rommem[20885] <= 16'hFFFF;
rommem[20886] <= 16'hFFFF;
rommem[20887] <= 16'hFFFF;
rommem[20888] <= 16'hFFFF;
rommem[20889] <= 16'hFFFF;
rommem[20890] <= 16'hFFFF;
rommem[20891] <= 16'hFFFF;
rommem[20892] <= 16'hFFFF;
rommem[20893] <= 16'hFFFF;
rommem[20894] <= 16'hFFFF;
rommem[20895] <= 16'hFFFF;
rommem[20896] <= 16'hFFFF;
rommem[20897] <= 16'hFFFF;
rommem[20898] <= 16'hFFFF;
rommem[20899] <= 16'hFFFF;
rommem[20900] <= 16'hFFFF;
rommem[20901] <= 16'hFFFF;
rommem[20902] <= 16'hFFFF;
rommem[20903] <= 16'hFFFF;
rommem[20904] <= 16'hFFFF;
rommem[20905] <= 16'hFFFF;
rommem[20906] <= 16'hFFFF;
rommem[20907] <= 16'hFFFF;
rommem[20908] <= 16'hFFFF;
rommem[20909] <= 16'hFFFF;
rommem[20910] <= 16'hFFFF;
rommem[20911] <= 16'hFFFF;
rommem[20912] <= 16'hFFFF;
rommem[20913] <= 16'hFFFF;
rommem[20914] <= 16'hFFFF;
rommem[20915] <= 16'hFFFF;
rommem[20916] <= 16'hFFFF;
rommem[20917] <= 16'hFFFF;
rommem[20918] <= 16'hFFFF;
rommem[20919] <= 16'hFFFF;
rommem[20920] <= 16'hFFFF;
rommem[20921] <= 16'hFFFF;
rommem[20922] <= 16'hFFFF;
rommem[20923] <= 16'hFFFF;
rommem[20924] <= 16'hFFFF;
rommem[20925] <= 16'hFFFF;
rommem[20926] <= 16'hFFFF;
rommem[20927] <= 16'hFFFF;
rommem[20928] <= 16'hFFFF;
rommem[20929] <= 16'hFFFF;
rommem[20930] <= 16'hFFFF;
rommem[20931] <= 16'hFFFF;
rommem[20932] <= 16'hFFFF;
rommem[20933] <= 16'hFFFF;
rommem[20934] <= 16'hFFFF;
rommem[20935] <= 16'hFFFF;
rommem[20936] <= 16'hFFFF;
rommem[20937] <= 16'hFFFF;
rommem[20938] <= 16'hFFFF;
rommem[20939] <= 16'hFFFF;
rommem[20940] <= 16'hFFFF;
rommem[20941] <= 16'hFFFF;
rommem[20942] <= 16'hFFFF;
rommem[20943] <= 16'hFFFF;
rommem[20944] <= 16'hFFFF;
rommem[20945] <= 16'hFFFF;
rommem[20946] <= 16'hFFFF;
rommem[20947] <= 16'hFFFF;
rommem[20948] <= 16'hFFFF;
rommem[20949] <= 16'hFFFF;
rommem[20950] <= 16'hFFFF;
rommem[20951] <= 16'hFFFF;
rommem[20952] <= 16'hFFFF;
rommem[20953] <= 16'hFFFF;
rommem[20954] <= 16'hFFFF;
rommem[20955] <= 16'hFFFF;
rommem[20956] <= 16'hFFFF;
rommem[20957] <= 16'hFFFF;
rommem[20958] <= 16'hFFFF;
rommem[20959] <= 16'hFFFF;
rommem[20960] <= 16'hFFFF;
rommem[20961] <= 16'hFFFF;
rommem[20962] <= 16'hFFFF;
rommem[20963] <= 16'hFFFF;
rommem[20964] <= 16'hFFFF;
rommem[20965] <= 16'hFFFF;
rommem[20966] <= 16'hFFFF;
rommem[20967] <= 16'hFFFF;
rommem[20968] <= 16'hFFFF;
rommem[20969] <= 16'hFFFF;
rommem[20970] <= 16'hFFFF;
rommem[20971] <= 16'hFFFF;
rommem[20972] <= 16'hFFFF;
rommem[20973] <= 16'hFFFF;
rommem[20974] <= 16'hFFFF;
rommem[20975] <= 16'hFFFF;
rommem[20976] <= 16'hFFFF;
rommem[20977] <= 16'hFFFF;
rommem[20978] <= 16'hFFFF;
rommem[20979] <= 16'hFFFF;
rommem[20980] <= 16'hFFFF;
rommem[20981] <= 16'hFFFF;
rommem[20982] <= 16'hFFFF;
rommem[20983] <= 16'hFFFF;
rommem[20984] <= 16'hFFFF;
rommem[20985] <= 16'hFFFF;
rommem[20986] <= 16'hFFFF;
rommem[20987] <= 16'hFFFF;
rommem[20988] <= 16'hFFFF;
rommem[20989] <= 16'hFFFF;
rommem[20990] <= 16'hFFFF;
rommem[20991] <= 16'hFFFF;
rommem[20992] <= 16'hFFFF;
rommem[20993] <= 16'hFFFF;
rommem[20994] <= 16'hFFFF;
rommem[20995] <= 16'hFFFF;
rommem[20996] <= 16'hFFFF;
rommem[20997] <= 16'hFFFF;
rommem[20998] <= 16'hFFFF;
rommem[20999] <= 16'hFFFF;
rommem[21000] <= 16'hFFFF;
rommem[21001] <= 16'hFFFF;
rommem[21002] <= 16'hFFFF;
rommem[21003] <= 16'hFFFF;
rommem[21004] <= 16'hFFFF;
rommem[21005] <= 16'hFFFF;
rommem[21006] <= 16'hFFFF;
rommem[21007] <= 16'hFFFF;
rommem[21008] <= 16'hFFFF;
rommem[21009] <= 16'hFFFF;
rommem[21010] <= 16'hFFFF;
rommem[21011] <= 16'hFFFF;
rommem[21012] <= 16'hFFFF;
rommem[21013] <= 16'hFFFF;
rommem[21014] <= 16'hFFFF;
rommem[21015] <= 16'hFFFF;
rommem[21016] <= 16'hFFFF;
rommem[21017] <= 16'hFFFF;
rommem[21018] <= 16'hFFFF;
rommem[21019] <= 16'hFFFF;
rommem[21020] <= 16'hFFFF;
rommem[21021] <= 16'hFFFF;
rommem[21022] <= 16'hFFFF;
rommem[21023] <= 16'hFFFF;
rommem[21024] <= 16'hFFFF;
rommem[21025] <= 16'hFFFF;
rommem[21026] <= 16'hFFFF;
rommem[21027] <= 16'hFFFF;
rommem[21028] <= 16'hFFFF;
rommem[21029] <= 16'hFFFF;
rommem[21030] <= 16'hFFFF;
rommem[21031] <= 16'hFFFF;
rommem[21032] <= 16'hFFFF;
rommem[21033] <= 16'hFFFF;
rommem[21034] <= 16'hFFFF;
rommem[21035] <= 16'hFFFF;
rommem[21036] <= 16'hFFFF;
rommem[21037] <= 16'hFFFF;
rommem[21038] <= 16'hFFFF;
rommem[21039] <= 16'hFFFF;
rommem[21040] <= 16'hFFFF;
rommem[21041] <= 16'hFFFF;
rommem[21042] <= 16'hFFFF;
rommem[21043] <= 16'hFFFF;
rommem[21044] <= 16'hFFFF;
rommem[21045] <= 16'hFFFF;
rommem[21046] <= 16'hFFFF;
rommem[21047] <= 16'hFFFF;
rommem[21048] <= 16'hFFFF;
rommem[21049] <= 16'hFFFF;
rommem[21050] <= 16'hFFFF;
rommem[21051] <= 16'hFFFF;
rommem[21052] <= 16'hFFFF;
rommem[21053] <= 16'hFFFF;
rommem[21054] <= 16'hFFFF;
rommem[21055] <= 16'hFFFF;
rommem[21056] <= 16'hFFFF;
rommem[21057] <= 16'hFFFF;
rommem[21058] <= 16'hFFFF;
rommem[21059] <= 16'hFFFF;
rommem[21060] <= 16'hFFFF;
rommem[21061] <= 16'hFFFF;
rommem[21062] <= 16'hFFFF;
rommem[21063] <= 16'hFFFF;
rommem[21064] <= 16'hFFFF;
rommem[21065] <= 16'hFFFF;
rommem[21066] <= 16'hFFFF;
rommem[21067] <= 16'hFFFF;
rommem[21068] <= 16'hFFFF;
rommem[21069] <= 16'hFFFF;
rommem[21070] <= 16'hFFFF;
rommem[21071] <= 16'hFFFF;
rommem[21072] <= 16'hFFFF;
rommem[21073] <= 16'hFFFF;
rommem[21074] <= 16'hFFFF;
rommem[21075] <= 16'hFFFF;
rommem[21076] <= 16'hFFFF;
rommem[21077] <= 16'hFFFF;
rommem[21078] <= 16'hFFFF;
rommem[21079] <= 16'hFFFF;
rommem[21080] <= 16'hFFFF;
rommem[21081] <= 16'hFFFF;
rommem[21082] <= 16'hFFFF;
rommem[21083] <= 16'hFFFF;
rommem[21084] <= 16'hFFFF;
rommem[21085] <= 16'hFFFF;
rommem[21086] <= 16'hFFFF;
rommem[21087] <= 16'hFFFF;
rommem[21088] <= 16'hFFFF;
rommem[21089] <= 16'hFFFF;
rommem[21090] <= 16'hFFFF;
rommem[21091] <= 16'hFFFF;
rommem[21092] <= 16'hFFFF;
rommem[21093] <= 16'hFFFF;
rommem[21094] <= 16'hFFFF;
rommem[21095] <= 16'hFFFF;
rommem[21096] <= 16'hFFFF;
rommem[21097] <= 16'hFFFF;
rommem[21098] <= 16'hFFFF;
rommem[21099] <= 16'hFFFF;
rommem[21100] <= 16'hFFFF;
rommem[21101] <= 16'hFFFF;
rommem[21102] <= 16'hFFFF;
rommem[21103] <= 16'hFFFF;
rommem[21104] <= 16'hFFFF;
rommem[21105] <= 16'hFFFF;
rommem[21106] <= 16'hFFFF;
rommem[21107] <= 16'hFFFF;
rommem[21108] <= 16'hFFFF;
rommem[21109] <= 16'hFFFF;
rommem[21110] <= 16'hFFFF;
rommem[21111] <= 16'hFFFF;
rommem[21112] <= 16'hFFFF;
rommem[21113] <= 16'hFFFF;
rommem[21114] <= 16'hFFFF;
rommem[21115] <= 16'hFFFF;
rommem[21116] <= 16'hFFFF;
rommem[21117] <= 16'hFFFF;
rommem[21118] <= 16'hFFFF;
rommem[21119] <= 16'hFFFF;
rommem[21120] <= 16'hFFFF;
rommem[21121] <= 16'hFFFF;
rommem[21122] <= 16'hFFFF;
rommem[21123] <= 16'hFFFF;
rommem[21124] <= 16'hFFFF;
rommem[21125] <= 16'hFFFF;
rommem[21126] <= 16'hFFFF;
rommem[21127] <= 16'hFFFF;
rommem[21128] <= 16'hFFFF;
rommem[21129] <= 16'hFFFF;
rommem[21130] <= 16'hFFFF;
rommem[21131] <= 16'hFFFF;
rommem[21132] <= 16'hFFFF;
rommem[21133] <= 16'hFFFF;
rommem[21134] <= 16'hFFFF;
rommem[21135] <= 16'hFFFF;
rommem[21136] <= 16'hFFFF;
rommem[21137] <= 16'hFFFF;
rommem[21138] <= 16'hFFFF;
rommem[21139] <= 16'hFFFF;
rommem[21140] <= 16'hFFFF;
rommem[21141] <= 16'hFFFF;
rommem[21142] <= 16'hFFFF;
rommem[21143] <= 16'hFFFF;
rommem[21144] <= 16'hFFFF;
rommem[21145] <= 16'hFFFF;
rommem[21146] <= 16'hFFFF;
rommem[21147] <= 16'hFFFF;
rommem[21148] <= 16'hFFFF;
rommem[21149] <= 16'hFFFF;
rommem[21150] <= 16'hFFFF;
rommem[21151] <= 16'hFFFF;
rommem[21152] <= 16'hFFFF;
rommem[21153] <= 16'hFFFF;
rommem[21154] <= 16'hFFFF;
rommem[21155] <= 16'hFFFF;
rommem[21156] <= 16'hFFFF;
rommem[21157] <= 16'hFFFF;
rommem[21158] <= 16'hFFFF;
rommem[21159] <= 16'hFFFF;
rommem[21160] <= 16'hFFFF;
rommem[21161] <= 16'hFFFF;
rommem[21162] <= 16'hFFFF;
rommem[21163] <= 16'hFFFF;
rommem[21164] <= 16'hFFFF;
rommem[21165] <= 16'hFFFF;
rommem[21166] <= 16'hFFFF;
rommem[21167] <= 16'hFFFF;
rommem[21168] <= 16'hFFFF;
rommem[21169] <= 16'hFFFF;
rommem[21170] <= 16'hFFFF;
rommem[21171] <= 16'hFFFF;
rommem[21172] <= 16'hFFFF;
rommem[21173] <= 16'hFFFF;
rommem[21174] <= 16'hFFFF;
rommem[21175] <= 16'hFFFF;
rommem[21176] <= 16'hFFFF;
rommem[21177] <= 16'hFFFF;
rommem[21178] <= 16'hFFFF;
rommem[21179] <= 16'hFFFF;
rommem[21180] <= 16'hFFFF;
rommem[21181] <= 16'hFFFF;
rommem[21182] <= 16'hFFFF;
rommem[21183] <= 16'hFFFF;
rommem[21184] <= 16'hFFFF;
rommem[21185] <= 16'hFFFF;
rommem[21186] <= 16'hFFFF;
rommem[21187] <= 16'hFFFF;
rommem[21188] <= 16'hFFFF;
rommem[21189] <= 16'hFFFF;
rommem[21190] <= 16'hFFFF;
rommem[21191] <= 16'hFFFF;
rommem[21192] <= 16'hFFFF;
rommem[21193] <= 16'hFFFF;
rommem[21194] <= 16'hFFFF;
rommem[21195] <= 16'hFFFF;
rommem[21196] <= 16'hFFFF;
rommem[21197] <= 16'hFFFF;
rommem[21198] <= 16'hFFFF;
rommem[21199] <= 16'hFFFF;
rommem[21200] <= 16'hFFFF;
rommem[21201] <= 16'hFFFF;
rommem[21202] <= 16'hFFFF;
rommem[21203] <= 16'hFFFF;
rommem[21204] <= 16'hFFFF;
rommem[21205] <= 16'hFFFF;
rommem[21206] <= 16'hFFFF;
rommem[21207] <= 16'hFFFF;
rommem[21208] <= 16'hFFFF;
rommem[21209] <= 16'hFFFF;
rommem[21210] <= 16'hFFFF;
rommem[21211] <= 16'hFFFF;
rommem[21212] <= 16'hFFFF;
rommem[21213] <= 16'hFFFF;
rommem[21214] <= 16'hFFFF;
rommem[21215] <= 16'hFFFF;
rommem[21216] <= 16'hFFFF;
rommem[21217] <= 16'hFFFF;
rommem[21218] <= 16'hFFFF;
rommem[21219] <= 16'hFFFF;
rommem[21220] <= 16'hFFFF;
rommem[21221] <= 16'hFFFF;
rommem[21222] <= 16'hFFFF;
rommem[21223] <= 16'hFFFF;
rommem[21224] <= 16'hFFFF;
rommem[21225] <= 16'hFFFF;
rommem[21226] <= 16'hFFFF;
rommem[21227] <= 16'hFFFF;
rommem[21228] <= 16'hFFFF;
rommem[21229] <= 16'hFFFF;
rommem[21230] <= 16'hFFFF;
rommem[21231] <= 16'hFFFF;
rommem[21232] <= 16'hFFFF;
rommem[21233] <= 16'hFFFF;
rommem[21234] <= 16'hFFFF;
rommem[21235] <= 16'hFFFF;
rommem[21236] <= 16'hFFFF;
rommem[21237] <= 16'hFFFF;
rommem[21238] <= 16'hFFFF;
rommem[21239] <= 16'hFFFF;
rommem[21240] <= 16'hFFFF;
rommem[21241] <= 16'hFFFF;
rommem[21242] <= 16'hFFFF;
rommem[21243] <= 16'hFFFF;
rommem[21244] <= 16'hFFFF;
rommem[21245] <= 16'hFFFF;
rommem[21246] <= 16'hFFFF;
rommem[21247] <= 16'hFFFF;
rommem[21248] <= 16'hFFFF;
rommem[21249] <= 16'hFFFF;
rommem[21250] <= 16'hFFFF;
rommem[21251] <= 16'hFFFF;
rommem[21252] <= 16'hFFFF;
rommem[21253] <= 16'hFFFF;
rommem[21254] <= 16'hFFFF;
rommem[21255] <= 16'hFFFF;
rommem[21256] <= 16'hFFFF;
rommem[21257] <= 16'hFFFF;
rommem[21258] <= 16'hFFFF;
rommem[21259] <= 16'hFFFF;
rommem[21260] <= 16'hFFFF;
rommem[21261] <= 16'hFFFF;
rommem[21262] <= 16'hFFFF;
rommem[21263] <= 16'hFFFF;
rommem[21264] <= 16'hFFFF;
rommem[21265] <= 16'hFFFF;
rommem[21266] <= 16'hFFFF;
rommem[21267] <= 16'hFFFF;
rommem[21268] <= 16'hFFFF;
rommem[21269] <= 16'hFFFF;
rommem[21270] <= 16'hFFFF;
rommem[21271] <= 16'hFFFF;
rommem[21272] <= 16'hFFFF;
rommem[21273] <= 16'hFFFF;
rommem[21274] <= 16'hFFFF;
rommem[21275] <= 16'hFFFF;
rommem[21276] <= 16'hFFFF;
rommem[21277] <= 16'hFFFF;
rommem[21278] <= 16'hFFFF;
rommem[21279] <= 16'hFFFF;
rommem[21280] <= 16'hFFFF;
rommem[21281] <= 16'hFFFF;
rommem[21282] <= 16'hFFFF;
rommem[21283] <= 16'hFFFF;
rommem[21284] <= 16'hFFFF;
rommem[21285] <= 16'hFFFF;
rommem[21286] <= 16'hFFFF;
rommem[21287] <= 16'hFFFF;
rommem[21288] <= 16'hFFFF;
rommem[21289] <= 16'hFFFF;
rommem[21290] <= 16'hFFFF;
rommem[21291] <= 16'hFFFF;
rommem[21292] <= 16'hFFFF;
rommem[21293] <= 16'hFFFF;
rommem[21294] <= 16'hFFFF;
rommem[21295] <= 16'hFFFF;
rommem[21296] <= 16'hFFFF;
rommem[21297] <= 16'hFFFF;
rommem[21298] <= 16'hFFFF;
rommem[21299] <= 16'hFFFF;
rommem[21300] <= 16'hFFFF;
rommem[21301] <= 16'hFFFF;
rommem[21302] <= 16'hFFFF;
rommem[21303] <= 16'hFFFF;
rommem[21304] <= 16'hFFFF;
rommem[21305] <= 16'hFFFF;
rommem[21306] <= 16'hFFFF;
rommem[21307] <= 16'hFFFF;
rommem[21308] <= 16'hFFFF;
rommem[21309] <= 16'hFFFF;
rommem[21310] <= 16'hFFFF;
rommem[21311] <= 16'hFFFF;
rommem[21312] <= 16'hFFFF;
rommem[21313] <= 16'hFFFF;
rommem[21314] <= 16'hFFFF;
rommem[21315] <= 16'hFFFF;
rommem[21316] <= 16'hFFFF;
rommem[21317] <= 16'hFFFF;
rommem[21318] <= 16'hFFFF;
rommem[21319] <= 16'hFFFF;
rommem[21320] <= 16'hFFFF;
rommem[21321] <= 16'hFFFF;
rommem[21322] <= 16'hFFFF;
rommem[21323] <= 16'hFFFF;
rommem[21324] <= 16'hFFFF;
rommem[21325] <= 16'hFFFF;
rommem[21326] <= 16'hFFFF;
rommem[21327] <= 16'hFFFF;
rommem[21328] <= 16'hFFFF;
rommem[21329] <= 16'hFFFF;
rommem[21330] <= 16'hFFFF;
rommem[21331] <= 16'hFFFF;
rommem[21332] <= 16'hFFFF;
rommem[21333] <= 16'hFFFF;
rommem[21334] <= 16'hFFFF;
rommem[21335] <= 16'hFFFF;
rommem[21336] <= 16'hFFFF;
rommem[21337] <= 16'hFFFF;
rommem[21338] <= 16'hFFFF;
rommem[21339] <= 16'hFFFF;
rommem[21340] <= 16'hFFFF;
rommem[21341] <= 16'hFFFF;
rommem[21342] <= 16'hFFFF;
rommem[21343] <= 16'hFFFF;
rommem[21344] <= 16'hFFFF;
rommem[21345] <= 16'hFFFF;
rommem[21346] <= 16'hFFFF;
rommem[21347] <= 16'hFFFF;
rommem[21348] <= 16'hFFFF;
rommem[21349] <= 16'hFFFF;
rommem[21350] <= 16'hFFFF;
rommem[21351] <= 16'hFFFF;
rommem[21352] <= 16'hFFFF;
rommem[21353] <= 16'hFFFF;
rommem[21354] <= 16'hFFFF;
rommem[21355] <= 16'hFFFF;
rommem[21356] <= 16'hFFFF;
rommem[21357] <= 16'hFFFF;
rommem[21358] <= 16'hFFFF;
rommem[21359] <= 16'hFFFF;
rommem[21360] <= 16'hFFFF;
rommem[21361] <= 16'hFFFF;
rommem[21362] <= 16'hFFFF;
rommem[21363] <= 16'hFFFF;
rommem[21364] <= 16'hFFFF;
rommem[21365] <= 16'hFFFF;
rommem[21366] <= 16'hFFFF;
rommem[21367] <= 16'hFFFF;
rommem[21368] <= 16'hFFFF;
rommem[21369] <= 16'hFFFF;
rommem[21370] <= 16'hFFFF;
rommem[21371] <= 16'hFFFF;
rommem[21372] <= 16'hFFFF;
rommem[21373] <= 16'hFFFF;
rommem[21374] <= 16'hFFFF;
rommem[21375] <= 16'hFFFF;
rommem[21376] <= 16'hFFFF;
rommem[21377] <= 16'hFFFF;
rommem[21378] <= 16'hFFFF;
rommem[21379] <= 16'hFFFF;
rommem[21380] <= 16'hFFFF;
rommem[21381] <= 16'hFFFF;
rommem[21382] <= 16'hFFFF;
rommem[21383] <= 16'hFFFF;
rommem[21384] <= 16'hFFFF;
rommem[21385] <= 16'hFFFF;
rommem[21386] <= 16'hFFFF;
rommem[21387] <= 16'hFFFF;
rommem[21388] <= 16'hFFFF;
rommem[21389] <= 16'hFFFF;
rommem[21390] <= 16'hFFFF;
rommem[21391] <= 16'hFFFF;
rommem[21392] <= 16'hFFFF;
rommem[21393] <= 16'hFFFF;
rommem[21394] <= 16'hFFFF;
rommem[21395] <= 16'hFFFF;
rommem[21396] <= 16'hFFFF;
rommem[21397] <= 16'hFFFF;
rommem[21398] <= 16'hFFFF;
rommem[21399] <= 16'hFFFF;
rommem[21400] <= 16'hFFFF;
rommem[21401] <= 16'hFFFF;
rommem[21402] <= 16'hFFFF;
rommem[21403] <= 16'hFFFF;
rommem[21404] <= 16'hFFFF;
rommem[21405] <= 16'hFFFF;
rommem[21406] <= 16'hFFFF;
rommem[21407] <= 16'hFFFF;
rommem[21408] <= 16'hFFFF;
rommem[21409] <= 16'hFFFF;
rommem[21410] <= 16'hFFFF;
rommem[21411] <= 16'hFFFF;
rommem[21412] <= 16'hFFFF;
rommem[21413] <= 16'hFFFF;
rommem[21414] <= 16'hFFFF;
rommem[21415] <= 16'hFFFF;
rommem[21416] <= 16'hFFFF;
rommem[21417] <= 16'hFFFF;
rommem[21418] <= 16'hFFFF;
rommem[21419] <= 16'hFFFF;
rommem[21420] <= 16'hFFFF;
rommem[21421] <= 16'hFFFF;
rommem[21422] <= 16'hFFFF;
rommem[21423] <= 16'hFFFF;
rommem[21424] <= 16'hFFFF;
rommem[21425] <= 16'hFFFF;
rommem[21426] <= 16'hFFFF;
rommem[21427] <= 16'hFFFF;
rommem[21428] <= 16'hFFFF;
rommem[21429] <= 16'hFFFF;
rommem[21430] <= 16'hFFFF;
rommem[21431] <= 16'hFFFF;
rommem[21432] <= 16'hFFFF;
rommem[21433] <= 16'hFFFF;
rommem[21434] <= 16'hFFFF;
rommem[21435] <= 16'hFFFF;
rommem[21436] <= 16'hFFFF;
rommem[21437] <= 16'hFFFF;
rommem[21438] <= 16'hFFFF;
rommem[21439] <= 16'hFFFF;
rommem[21440] <= 16'hFFFF;
rommem[21441] <= 16'hFFFF;
rommem[21442] <= 16'hFFFF;
rommem[21443] <= 16'hFFFF;
rommem[21444] <= 16'hFFFF;
rommem[21445] <= 16'hFFFF;
rommem[21446] <= 16'hFFFF;
rommem[21447] <= 16'hFFFF;
rommem[21448] <= 16'hFFFF;
rommem[21449] <= 16'hFFFF;
rommem[21450] <= 16'hFFFF;
rommem[21451] <= 16'hFFFF;
rommem[21452] <= 16'hFFFF;
rommem[21453] <= 16'hFFFF;
rommem[21454] <= 16'hFFFF;
rommem[21455] <= 16'hFFFF;
rommem[21456] <= 16'hFFFF;
rommem[21457] <= 16'hFFFF;
rommem[21458] <= 16'hFFFF;
rommem[21459] <= 16'hFFFF;
rommem[21460] <= 16'hFFFF;
rommem[21461] <= 16'hFFFF;
rommem[21462] <= 16'hFFFF;
rommem[21463] <= 16'hFFFF;
rommem[21464] <= 16'hFFFF;
rommem[21465] <= 16'hFFFF;
rommem[21466] <= 16'hFFFF;
rommem[21467] <= 16'hFFFF;
rommem[21468] <= 16'hFFFF;
rommem[21469] <= 16'hFFFF;
rommem[21470] <= 16'hFFFF;
rommem[21471] <= 16'hFFFF;
rommem[21472] <= 16'hFFFF;
rommem[21473] <= 16'hFFFF;
rommem[21474] <= 16'hFFFF;
rommem[21475] <= 16'hFFFF;
rommem[21476] <= 16'hFFFF;
rommem[21477] <= 16'hFFFF;
rommem[21478] <= 16'hFFFF;
rommem[21479] <= 16'hFFFF;
rommem[21480] <= 16'hFFFF;
rommem[21481] <= 16'hFFFF;
rommem[21482] <= 16'hFFFF;
rommem[21483] <= 16'hFFFF;
rommem[21484] <= 16'hFFFF;
rommem[21485] <= 16'hFFFF;
rommem[21486] <= 16'hFFFF;
rommem[21487] <= 16'hFFFF;
rommem[21488] <= 16'hFFFF;
rommem[21489] <= 16'hFFFF;
rommem[21490] <= 16'hFFFF;
rommem[21491] <= 16'hFFFF;
rommem[21492] <= 16'hFFFF;
rommem[21493] <= 16'hFFFF;
rommem[21494] <= 16'hFFFF;
rommem[21495] <= 16'hFFFF;
rommem[21496] <= 16'hFFFF;
rommem[21497] <= 16'hFFFF;
rommem[21498] <= 16'hFFFF;
rommem[21499] <= 16'hFFFF;
rommem[21500] <= 16'hFFFF;
rommem[21501] <= 16'hFFFF;
rommem[21502] <= 16'hFFFF;
rommem[21503] <= 16'hFFFF;
rommem[21504] <= 16'hFFFF;
rommem[21505] <= 16'hFFFF;
rommem[21506] <= 16'hFFFF;
rommem[21507] <= 16'hFFFF;
rommem[21508] <= 16'hFFFF;
rommem[21509] <= 16'hFFFF;
rommem[21510] <= 16'hFFFF;
rommem[21511] <= 16'hFFFF;
rommem[21512] <= 16'hFFFF;
rommem[21513] <= 16'hFFFF;
rommem[21514] <= 16'hFFFF;
rommem[21515] <= 16'hFFFF;
rommem[21516] <= 16'hFFFF;
rommem[21517] <= 16'hFFFF;
rommem[21518] <= 16'hFFFF;
rommem[21519] <= 16'hFFFF;
rommem[21520] <= 16'hFFFF;
rommem[21521] <= 16'hFFFF;
rommem[21522] <= 16'hFFFF;
rommem[21523] <= 16'hFFFF;
rommem[21524] <= 16'hFFFF;
rommem[21525] <= 16'hFFFF;
rommem[21526] <= 16'hFFFF;
rommem[21527] <= 16'hFFFF;
rommem[21528] <= 16'hFFFF;
rommem[21529] <= 16'hFFFF;
rommem[21530] <= 16'hFFFF;
rommem[21531] <= 16'hFFFF;
rommem[21532] <= 16'hFFFF;
rommem[21533] <= 16'hFFFF;
rommem[21534] <= 16'hFFFF;
rommem[21535] <= 16'hFFFF;
rommem[21536] <= 16'hFFFF;
rommem[21537] <= 16'hFFFF;
rommem[21538] <= 16'hFFFF;
rommem[21539] <= 16'hFFFF;
rommem[21540] <= 16'hFFFF;
rommem[21541] <= 16'hFFFF;
rommem[21542] <= 16'hFFFF;
rommem[21543] <= 16'hFFFF;
rommem[21544] <= 16'hFFFF;
rommem[21545] <= 16'hFFFF;
rommem[21546] <= 16'hFFFF;
rommem[21547] <= 16'hFFFF;
rommem[21548] <= 16'hFFFF;
rommem[21549] <= 16'hFFFF;
rommem[21550] <= 16'hFFFF;
rommem[21551] <= 16'hFFFF;
rommem[21552] <= 16'hFFFF;
rommem[21553] <= 16'hFFFF;
rommem[21554] <= 16'hFFFF;
rommem[21555] <= 16'hFFFF;
rommem[21556] <= 16'hFFFF;
rommem[21557] <= 16'hFFFF;
rommem[21558] <= 16'hFFFF;
rommem[21559] <= 16'hFFFF;
rommem[21560] <= 16'hFFFF;
rommem[21561] <= 16'hFFFF;
rommem[21562] <= 16'hFFFF;
rommem[21563] <= 16'hFFFF;
rommem[21564] <= 16'hFFFF;
rommem[21565] <= 16'hFFFF;
rommem[21566] <= 16'hFFFF;
rommem[21567] <= 16'hFFFF;
rommem[21568] <= 16'hFFFF;
rommem[21569] <= 16'hFFFF;
rommem[21570] <= 16'hFFFF;
rommem[21571] <= 16'hFFFF;
rommem[21572] <= 16'hFFFF;
rommem[21573] <= 16'hFFFF;
rommem[21574] <= 16'hFFFF;
rommem[21575] <= 16'hFFFF;
rommem[21576] <= 16'hFFFF;
rommem[21577] <= 16'hFFFF;
rommem[21578] <= 16'hFFFF;
rommem[21579] <= 16'hFFFF;
rommem[21580] <= 16'hFFFF;
rommem[21581] <= 16'hFFFF;
rommem[21582] <= 16'hFFFF;
rommem[21583] <= 16'hFFFF;
rommem[21584] <= 16'hFFFF;
rommem[21585] <= 16'hFFFF;
rommem[21586] <= 16'hFFFF;
rommem[21587] <= 16'hFFFF;
rommem[21588] <= 16'hFFFF;
rommem[21589] <= 16'hFFFF;
rommem[21590] <= 16'hFFFF;
rommem[21591] <= 16'hFFFF;
rommem[21592] <= 16'hFFFF;
rommem[21593] <= 16'hFFFF;
rommem[21594] <= 16'hFFFF;
rommem[21595] <= 16'hFFFF;
rommem[21596] <= 16'hFFFF;
rommem[21597] <= 16'hFFFF;
rommem[21598] <= 16'hFFFF;
rommem[21599] <= 16'hFFFF;
rommem[21600] <= 16'hFFFF;
rommem[21601] <= 16'hFFFF;
rommem[21602] <= 16'hFFFF;
rommem[21603] <= 16'hFFFF;
rommem[21604] <= 16'hFFFF;
rommem[21605] <= 16'hFFFF;
rommem[21606] <= 16'hFFFF;
rommem[21607] <= 16'hFFFF;
rommem[21608] <= 16'hFFFF;
rommem[21609] <= 16'hFFFF;
rommem[21610] <= 16'hFFFF;
rommem[21611] <= 16'hFFFF;
rommem[21612] <= 16'hFFFF;
rommem[21613] <= 16'hFFFF;
rommem[21614] <= 16'hFFFF;
rommem[21615] <= 16'hFFFF;
rommem[21616] <= 16'hFFFF;
rommem[21617] <= 16'hFFFF;
rommem[21618] <= 16'hFFFF;
rommem[21619] <= 16'hFFFF;
rommem[21620] <= 16'hFFFF;
rommem[21621] <= 16'hFFFF;
rommem[21622] <= 16'hFFFF;
rommem[21623] <= 16'hFFFF;
rommem[21624] <= 16'hFFFF;
rommem[21625] <= 16'hFFFF;
rommem[21626] <= 16'hFFFF;
rommem[21627] <= 16'hFFFF;
rommem[21628] <= 16'hFFFF;
rommem[21629] <= 16'hFFFF;
rommem[21630] <= 16'hFFFF;
rommem[21631] <= 16'hFFFF;
rommem[21632] <= 16'hFFFF;
rommem[21633] <= 16'hFFFF;
rommem[21634] <= 16'hFFFF;
rommem[21635] <= 16'hFFFF;
rommem[21636] <= 16'hFFFF;
rommem[21637] <= 16'hFFFF;
rommem[21638] <= 16'hFFFF;
rommem[21639] <= 16'hFFFF;
rommem[21640] <= 16'hFFFF;
rommem[21641] <= 16'hFFFF;
rommem[21642] <= 16'hFFFF;
rommem[21643] <= 16'hFFFF;
rommem[21644] <= 16'hFFFF;
rommem[21645] <= 16'hFFFF;
rommem[21646] <= 16'hFFFF;
rommem[21647] <= 16'hFFFF;
rommem[21648] <= 16'hFFFF;
rommem[21649] <= 16'hFFFF;
rommem[21650] <= 16'hFFFF;
rommem[21651] <= 16'hFFFF;
rommem[21652] <= 16'hFFFF;
rommem[21653] <= 16'hFFFF;
rommem[21654] <= 16'hFFFF;
rommem[21655] <= 16'hFFFF;
rommem[21656] <= 16'hFFFF;
rommem[21657] <= 16'hFFFF;
rommem[21658] <= 16'hFFFF;
rommem[21659] <= 16'hFFFF;
rommem[21660] <= 16'hFFFF;
rommem[21661] <= 16'hFFFF;
rommem[21662] <= 16'hFFFF;
rommem[21663] <= 16'hFFFF;
rommem[21664] <= 16'hFFFF;
rommem[21665] <= 16'hFFFF;
rommem[21666] <= 16'hFFFF;
rommem[21667] <= 16'hFFFF;
rommem[21668] <= 16'hFFFF;
rommem[21669] <= 16'hFFFF;
rommem[21670] <= 16'hFFFF;
rommem[21671] <= 16'hFFFF;
rommem[21672] <= 16'hFFFF;
rommem[21673] <= 16'hFFFF;
rommem[21674] <= 16'hFFFF;
rommem[21675] <= 16'hFFFF;
rommem[21676] <= 16'hFFFF;
rommem[21677] <= 16'hFFFF;
rommem[21678] <= 16'hFFFF;
rommem[21679] <= 16'hFFFF;
rommem[21680] <= 16'hFFFF;
rommem[21681] <= 16'hFFFF;
rommem[21682] <= 16'hFFFF;
rommem[21683] <= 16'hFFFF;
rommem[21684] <= 16'hFFFF;
rommem[21685] <= 16'hFFFF;
rommem[21686] <= 16'hFFFF;
rommem[21687] <= 16'hFFFF;
rommem[21688] <= 16'hFFFF;
rommem[21689] <= 16'hFFFF;
rommem[21690] <= 16'hFFFF;
rommem[21691] <= 16'hFFFF;
rommem[21692] <= 16'hFFFF;
rommem[21693] <= 16'hFFFF;
rommem[21694] <= 16'hFFFF;
rommem[21695] <= 16'hFFFF;
rommem[21696] <= 16'hFFFF;
rommem[21697] <= 16'hFFFF;
rommem[21698] <= 16'hFFFF;
rommem[21699] <= 16'hFFFF;
rommem[21700] <= 16'hFFFF;
rommem[21701] <= 16'hFFFF;
rommem[21702] <= 16'hFFFF;
rommem[21703] <= 16'hFFFF;
rommem[21704] <= 16'hFFFF;
rommem[21705] <= 16'hFFFF;
rommem[21706] <= 16'hFFFF;
rommem[21707] <= 16'hFFFF;
rommem[21708] <= 16'hFFFF;
rommem[21709] <= 16'hFFFF;
rommem[21710] <= 16'hFFFF;
rommem[21711] <= 16'hFFFF;
rommem[21712] <= 16'hFFFF;
rommem[21713] <= 16'hFFFF;
rommem[21714] <= 16'hFFFF;
rommem[21715] <= 16'hFFFF;
rommem[21716] <= 16'hFFFF;
rommem[21717] <= 16'hFFFF;
rommem[21718] <= 16'hFFFF;
rommem[21719] <= 16'hFFFF;
rommem[21720] <= 16'hFFFF;
rommem[21721] <= 16'hFFFF;
rommem[21722] <= 16'hFFFF;
rommem[21723] <= 16'hFFFF;
rommem[21724] <= 16'hFFFF;
rommem[21725] <= 16'hFFFF;
rommem[21726] <= 16'hFFFF;
rommem[21727] <= 16'hFFFF;
rommem[21728] <= 16'hFFFF;
rommem[21729] <= 16'hFFFF;
rommem[21730] <= 16'hFFFF;
rommem[21731] <= 16'hFFFF;
rommem[21732] <= 16'hFFFF;
rommem[21733] <= 16'hFFFF;
rommem[21734] <= 16'hFFFF;
rommem[21735] <= 16'hFFFF;
rommem[21736] <= 16'hFFFF;
rommem[21737] <= 16'hFFFF;
rommem[21738] <= 16'hFFFF;
rommem[21739] <= 16'hFFFF;
rommem[21740] <= 16'hFFFF;
rommem[21741] <= 16'hFFFF;
rommem[21742] <= 16'hFFFF;
rommem[21743] <= 16'hFFFF;
rommem[21744] <= 16'hFFFF;
rommem[21745] <= 16'hFFFF;
rommem[21746] <= 16'hFFFF;
rommem[21747] <= 16'hFFFF;
rommem[21748] <= 16'hFFFF;
rommem[21749] <= 16'hFFFF;
rommem[21750] <= 16'hFFFF;
rommem[21751] <= 16'hFFFF;
rommem[21752] <= 16'hFFFF;
rommem[21753] <= 16'hFFFF;
rommem[21754] <= 16'hFFFF;
rommem[21755] <= 16'hFFFF;
rommem[21756] <= 16'hFFFF;
rommem[21757] <= 16'hFFFF;
rommem[21758] <= 16'hFFFF;
rommem[21759] <= 16'hFFFF;
rommem[21760] <= 16'hFFFF;
rommem[21761] <= 16'hFFFF;
rommem[21762] <= 16'hFFFF;
rommem[21763] <= 16'hFFFF;
rommem[21764] <= 16'hFFFF;
rommem[21765] <= 16'hFFFF;
rommem[21766] <= 16'hFFFF;
rommem[21767] <= 16'hFFFF;
rommem[21768] <= 16'hFFFF;
rommem[21769] <= 16'hFFFF;
rommem[21770] <= 16'hFFFF;
rommem[21771] <= 16'hFFFF;
rommem[21772] <= 16'hFFFF;
rommem[21773] <= 16'hFFFF;
rommem[21774] <= 16'hFFFF;
rommem[21775] <= 16'hFFFF;
rommem[21776] <= 16'hFFFF;
rommem[21777] <= 16'hFFFF;
rommem[21778] <= 16'hFFFF;
rommem[21779] <= 16'hFFFF;
rommem[21780] <= 16'hFFFF;
rommem[21781] <= 16'hFFFF;
rommem[21782] <= 16'hFFFF;
rommem[21783] <= 16'hFFFF;
rommem[21784] <= 16'hFFFF;
rommem[21785] <= 16'hFFFF;
rommem[21786] <= 16'hFFFF;
rommem[21787] <= 16'hFFFF;
rommem[21788] <= 16'hFFFF;
rommem[21789] <= 16'hFFFF;
rommem[21790] <= 16'hFFFF;
rommem[21791] <= 16'hFFFF;
rommem[21792] <= 16'hFFFF;
rommem[21793] <= 16'hFFFF;
rommem[21794] <= 16'hFFFF;
rommem[21795] <= 16'hFFFF;
rommem[21796] <= 16'hFFFF;
rommem[21797] <= 16'hFFFF;
rommem[21798] <= 16'hFFFF;
rommem[21799] <= 16'hFFFF;
rommem[21800] <= 16'hFFFF;
rommem[21801] <= 16'hFFFF;
rommem[21802] <= 16'hFFFF;
rommem[21803] <= 16'hFFFF;
rommem[21804] <= 16'hFFFF;
rommem[21805] <= 16'hFFFF;
rommem[21806] <= 16'hFFFF;
rommem[21807] <= 16'hFFFF;
rommem[21808] <= 16'hFFFF;
rommem[21809] <= 16'hFFFF;
rommem[21810] <= 16'hFFFF;
rommem[21811] <= 16'hFFFF;
rommem[21812] <= 16'hFFFF;
rommem[21813] <= 16'hFFFF;
rommem[21814] <= 16'hFFFF;
rommem[21815] <= 16'hFFFF;
rommem[21816] <= 16'hFFFF;
rommem[21817] <= 16'hFFFF;
rommem[21818] <= 16'hFFFF;
rommem[21819] <= 16'hFFFF;
rommem[21820] <= 16'hFFFF;
rommem[21821] <= 16'hFFFF;
rommem[21822] <= 16'hFFFF;
rommem[21823] <= 16'hFFFF;
rommem[21824] <= 16'hFFFF;
rommem[21825] <= 16'hFFFF;
rommem[21826] <= 16'hFFFF;
rommem[21827] <= 16'hFFFF;
rommem[21828] <= 16'hFFFF;
rommem[21829] <= 16'hFFFF;
rommem[21830] <= 16'hFFFF;
rommem[21831] <= 16'hFFFF;
rommem[21832] <= 16'hFFFF;
rommem[21833] <= 16'hFFFF;
rommem[21834] <= 16'hFFFF;
rommem[21835] <= 16'hFFFF;
rommem[21836] <= 16'hFFFF;
rommem[21837] <= 16'hFFFF;
rommem[21838] <= 16'hFFFF;
rommem[21839] <= 16'hFFFF;
rommem[21840] <= 16'hFFFF;
rommem[21841] <= 16'hFFFF;
rommem[21842] <= 16'hFFFF;
rommem[21843] <= 16'hFFFF;
rommem[21844] <= 16'hFFFF;
rommem[21845] <= 16'hFFFF;
rommem[21846] <= 16'hFFFF;
rommem[21847] <= 16'hFFFF;
rommem[21848] <= 16'hFFFF;
rommem[21849] <= 16'hFFFF;
rommem[21850] <= 16'hFFFF;
rommem[21851] <= 16'hFFFF;
rommem[21852] <= 16'hFFFF;
rommem[21853] <= 16'hFFFF;
rommem[21854] <= 16'hFFFF;
rommem[21855] <= 16'hFFFF;
rommem[21856] <= 16'hFFFF;
rommem[21857] <= 16'hFFFF;
rommem[21858] <= 16'hFFFF;
rommem[21859] <= 16'hFFFF;
rommem[21860] <= 16'hFFFF;
rommem[21861] <= 16'hFFFF;
rommem[21862] <= 16'hFFFF;
rommem[21863] <= 16'hFFFF;
rommem[21864] <= 16'hFFFF;
rommem[21865] <= 16'hFFFF;
rommem[21866] <= 16'hFFFF;
rommem[21867] <= 16'hFFFF;
rommem[21868] <= 16'hFFFF;
rommem[21869] <= 16'hFFFF;
rommem[21870] <= 16'hFFFF;
rommem[21871] <= 16'hFFFF;
rommem[21872] <= 16'hFFFF;
rommem[21873] <= 16'hFFFF;
rommem[21874] <= 16'hFFFF;
rommem[21875] <= 16'hFFFF;
rommem[21876] <= 16'hFFFF;
rommem[21877] <= 16'hFFFF;
rommem[21878] <= 16'hFFFF;
rommem[21879] <= 16'hFFFF;
rommem[21880] <= 16'hFFFF;
rommem[21881] <= 16'hFFFF;
rommem[21882] <= 16'hFFFF;
rommem[21883] <= 16'hFFFF;
rommem[21884] <= 16'hFFFF;
rommem[21885] <= 16'hFFFF;
rommem[21886] <= 16'hFFFF;
rommem[21887] <= 16'hFFFF;
rommem[21888] <= 16'hFFFF;
rommem[21889] <= 16'hFFFF;
rommem[21890] <= 16'hFFFF;
rommem[21891] <= 16'hFFFF;
rommem[21892] <= 16'hFFFF;
rommem[21893] <= 16'hFFFF;
rommem[21894] <= 16'hFFFF;
rommem[21895] <= 16'hFFFF;
rommem[21896] <= 16'hFFFF;
rommem[21897] <= 16'hFFFF;
rommem[21898] <= 16'hFFFF;
rommem[21899] <= 16'hFFFF;
rommem[21900] <= 16'hFFFF;
rommem[21901] <= 16'hFFFF;
rommem[21902] <= 16'hFFFF;
rommem[21903] <= 16'hFFFF;
rommem[21904] <= 16'hFFFF;
rommem[21905] <= 16'hFFFF;
rommem[21906] <= 16'hFFFF;
rommem[21907] <= 16'hFFFF;
rommem[21908] <= 16'hFFFF;
rommem[21909] <= 16'hFFFF;
rommem[21910] <= 16'hFFFF;
rommem[21911] <= 16'hFFFF;
rommem[21912] <= 16'hFFFF;
rommem[21913] <= 16'hFFFF;
rommem[21914] <= 16'hFFFF;
rommem[21915] <= 16'hFFFF;
rommem[21916] <= 16'hFFFF;
rommem[21917] <= 16'hFFFF;
rommem[21918] <= 16'hFFFF;
rommem[21919] <= 16'hFFFF;
rommem[21920] <= 16'hFFFF;
rommem[21921] <= 16'hFFFF;
rommem[21922] <= 16'hFFFF;
rommem[21923] <= 16'hFFFF;
rommem[21924] <= 16'hFFFF;
rommem[21925] <= 16'hFFFF;
rommem[21926] <= 16'hFFFF;
rommem[21927] <= 16'hFFFF;
rommem[21928] <= 16'hFFFF;
rommem[21929] <= 16'hFFFF;
rommem[21930] <= 16'hFFFF;
rommem[21931] <= 16'hFFFF;
rommem[21932] <= 16'hFFFF;
rommem[21933] <= 16'hFFFF;
rommem[21934] <= 16'hFFFF;
rommem[21935] <= 16'hFFFF;
rommem[21936] <= 16'hFFFF;
rommem[21937] <= 16'hFFFF;
rommem[21938] <= 16'hFFFF;
rommem[21939] <= 16'hFFFF;
rommem[21940] <= 16'hFFFF;
rommem[21941] <= 16'hFFFF;
rommem[21942] <= 16'hFFFF;
rommem[21943] <= 16'hFFFF;
rommem[21944] <= 16'hFFFF;
rommem[21945] <= 16'hFFFF;
rommem[21946] <= 16'hFFFF;
rommem[21947] <= 16'hFFFF;
rommem[21948] <= 16'hFFFF;
rommem[21949] <= 16'hFFFF;
rommem[21950] <= 16'hFFFF;
rommem[21951] <= 16'hFFFF;
rommem[21952] <= 16'hFFFF;
rommem[21953] <= 16'hFFFF;
rommem[21954] <= 16'hFFFF;
rommem[21955] <= 16'hFFFF;
rommem[21956] <= 16'hFFFF;
rommem[21957] <= 16'hFFFF;
rommem[21958] <= 16'hFFFF;
rommem[21959] <= 16'hFFFF;
rommem[21960] <= 16'hFFFF;
rommem[21961] <= 16'hFFFF;
rommem[21962] <= 16'hFFFF;
rommem[21963] <= 16'hFFFF;
rommem[21964] <= 16'hFFFF;
rommem[21965] <= 16'hFFFF;
rommem[21966] <= 16'hFFFF;
rommem[21967] <= 16'hFFFF;
rommem[21968] <= 16'hFFFF;
rommem[21969] <= 16'hFFFF;
rommem[21970] <= 16'hFFFF;
rommem[21971] <= 16'hFFFF;
rommem[21972] <= 16'hFFFF;
rommem[21973] <= 16'hFFFF;
rommem[21974] <= 16'hFFFF;
rommem[21975] <= 16'hFFFF;
rommem[21976] <= 16'hFFFF;
rommem[21977] <= 16'hFFFF;
rommem[21978] <= 16'hFFFF;
rommem[21979] <= 16'hFFFF;
rommem[21980] <= 16'hFFFF;
rommem[21981] <= 16'hFFFF;
rommem[21982] <= 16'hFFFF;
rommem[21983] <= 16'hFFFF;
rommem[21984] <= 16'hFFFF;
rommem[21985] <= 16'hFFFF;
rommem[21986] <= 16'hFFFF;
rommem[21987] <= 16'hFFFF;
rommem[21988] <= 16'hFFFF;
rommem[21989] <= 16'hFFFF;
rommem[21990] <= 16'hFFFF;
rommem[21991] <= 16'hFFFF;
rommem[21992] <= 16'hFFFF;
rommem[21993] <= 16'hFFFF;
rommem[21994] <= 16'hFFFF;
rommem[21995] <= 16'hFFFF;
rommem[21996] <= 16'hFFFF;
rommem[21997] <= 16'hFFFF;
rommem[21998] <= 16'hFFFF;
rommem[21999] <= 16'hFFFF;
rommem[22000] <= 16'hFFFF;
rommem[22001] <= 16'hFFFF;
rommem[22002] <= 16'hFFFF;
rommem[22003] <= 16'hFFFF;
rommem[22004] <= 16'hFFFF;
rommem[22005] <= 16'hFFFF;
rommem[22006] <= 16'hFFFF;
rommem[22007] <= 16'hFFFF;
rommem[22008] <= 16'hFFFF;
rommem[22009] <= 16'hFFFF;
rommem[22010] <= 16'hFFFF;
rommem[22011] <= 16'hFFFF;
rommem[22012] <= 16'hFFFF;
rommem[22013] <= 16'hFFFF;
rommem[22014] <= 16'hFFFF;
rommem[22015] <= 16'hFFFF;
rommem[22016] <= 16'hFFFF;
rommem[22017] <= 16'hFFFF;
rommem[22018] <= 16'hFFFF;
rommem[22019] <= 16'hFFFF;
rommem[22020] <= 16'hFFFF;
rommem[22021] <= 16'hFFFF;
rommem[22022] <= 16'hFFFF;
rommem[22023] <= 16'hFFFF;
rommem[22024] <= 16'hFFFF;
rommem[22025] <= 16'hFFFF;
rommem[22026] <= 16'hFFFF;
rommem[22027] <= 16'hFFFF;
rommem[22028] <= 16'hFFFF;
rommem[22029] <= 16'hFFFF;
rommem[22030] <= 16'hFFFF;
rommem[22031] <= 16'hFFFF;
rommem[22032] <= 16'hFFFF;
rommem[22033] <= 16'hFFFF;
rommem[22034] <= 16'hFFFF;
rommem[22035] <= 16'hFFFF;
rommem[22036] <= 16'hFFFF;
rommem[22037] <= 16'hFFFF;
rommem[22038] <= 16'hFFFF;
rommem[22039] <= 16'hFFFF;
rommem[22040] <= 16'hFFFF;
rommem[22041] <= 16'hFFFF;
rommem[22042] <= 16'hFFFF;
rommem[22043] <= 16'hFFFF;
rommem[22044] <= 16'hFFFF;
rommem[22045] <= 16'hFFFF;
rommem[22046] <= 16'hFFFF;
rommem[22047] <= 16'hFFFF;
rommem[22048] <= 16'hFFFF;
rommem[22049] <= 16'hFFFF;
rommem[22050] <= 16'hFFFF;
rommem[22051] <= 16'hFFFF;
rommem[22052] <= 16'hFFFF;
rommem[22053] <= 16'hFFFF;
rommem[22054] <= 16'hFFFF;
rommem[22055] <= 16'hFFFF;
rommem[22056] <= 16'hFFFF;
rommem[22057] <= 16'hFFFF;
rommem[22058] <= 16'hFFFF;
rommem[22059] <= 16'hFFFF;
rommem[22060] <= 16'hFFFF;
rommem[22061] <= 16'hFFFF;
rommem[22062] <= 16'hFFFF;
rommem[22063] <= 16'hFFFF;
rommem[22064] <= 16'hFFFF;
rommem[22065] <= 16'hFFFF;
rommem[22066] <= 16'hFFFF;
rommem[22067] <= 16'hFFFF;
rommem[22068] <= 16'hFFFF;
rommem[22069] <= 16'hFFFF;
rommem[22070] <= 16'hFFFF;
rommem[22071] <= 16'hFFFF;
rommem[22072] <= 16'hFFFF;
rommem[22073] <= 16'hFFFF;
rommem[22074] <= 16'hFFFF;
rommem[22075] <= 16'hFFFF;
rommem[22076] <= 16'hFFFF;
rommem[22077] <= 16'hFFFF;
rommem[22078] <= 16'hFFFF;
rommem[22079] <= 16'hFFFF;
rommem[22080] <= 16'hFFFF;
rommem[22081] <= 16'hFFFF;
rommem[22082] <= 16'hFFFF;
rommem[22083] <= 16'hFFFF;
rommem[22084] <= 16'hFFFF;
rommem[22085] <= 16'hFFFF;
rommem[22086] <= 16'hFFFF;
rommem[22087] <= 16'hFFFF;
rommem[22088] <= 16'hFFFF;
rommem[22089] <= 16'hFFFF;
rommem[22090] <= 16'hFFFF;
rommem[22091] <= 16'hFFFF;
rommem[22092] <= 16'hFFFF;
rommem[22093] <= 16'hFFFF;
rommem[22094] <= 16'hFFFF;
rommem[22095] <= 16'hFFFF;
rommem[22096] <= 16'hFFFF;
rommem[22097] <= 16'hFFFF;
rommem[22098] <= 16'hFFFF;
rommem[22099] <= 16'hFFFF;
rommem[22100] <= 16'hFFFF;
rommem[22101] <= 16'hFFFF;
rommem[22102] <= 16'hFFFF;
rommem[22103] <= 16'hFFFF;
rommem[22104] <= 16'hFFFF;
rommem[22105] <= 16'hFFFF;
rommem[22106] <= 16'hFFFF;
rommem[22107] <= 16'hFFFF;
rommem[22108] <= 16'hFFFF;
rommem[22109] <= 16'hFFFF;
rommem[22110] <= 16'hFFFF;
rommem[22111] <= 16'hFFFF;
rommem[22112] <= 16'hFFFF;
rommem[22113] <= 16'hFFFF;
rommem[22114] <= 16'hFFFF;
rommem[22115] <= 16'hFFFF;
rommem[22116] <= 16'hFFFF;
rommem[22117] <= 16'hFFFF;
rommem[22118] <= 16'hFFFF;
rommem[22119] <= 16'hFFFF;
rommem[22120] <= 16'hFFFF;
rommem[22121] <= 16'hFFFF;
rommem[22122] <= 16'hFFFF;
rommem[22123] <= 16'hFFFF;
rommem[22124] <= 16'hFFFF;
rommem[22125] <= 16'hFFFF;
rommem[22126] <= 16'hFFFF;
rommem[22127] <= 16'hFFFF;
rommem[22128] <= 16'hFFFF;
rommem[22129] <= 16'hFFFF;
rommem[22130] <= 16'hFFFF;
rommem[22131] <= 16'hFFFF;
rommem[22132] <= 16'hFFFF;
rommem[22133] <= 16'hFFFF;
rommem[22134] <= 16'hFFFF;
rommem[22135] <= 16'hFFFF;
rommem[22136] <= 16'hFFFF;
rommem[22137] <= 16'hFFFF;
rommem[22138] <= 16'hFFFF;
rommem[22139] <= 16'hFFFF;
rommem[22140] <= 16'hFFFF;
rommem[22141] <= 16'hFFFF;
rommem[22142] <= 16'hFFFF;
rommem[22143] <= 16'hFFFF;
rommem[22144] <= 16'hFFFF;
rommem[22145] <= 16'hFFFF;
rommem[22146] <= 16'hFFFF;
rommem[22147] <= 16'hFFFF;
rommem[22148] <= 16'hFFFF;
rommem[22149] <= 16'hFFFF;
rommem[22150] <= 16'hFFFF;
rommem[22151] <= 16'hFFFF;
rommem[22152] <= 16'hFFFF;
rommem[22153] <= 16'hFFFF;
rommem[22154] <= 16'hFFFF;
rommem[22155] <= 16'hFFFF;
rommem[22156] <= 16'hFFFF;
rommem[22157] <= 16'hFFFF;
rommem[22158] <= 16'hFFFF;
rommem[22159] <= 16'hFFFF;
rommem[22160] <= 16'hFFFF;
rommem[22161] <= 16'hFFFF;
rommem[22162] <= 16'hFFFF;
rommem[22163] <= 16'hFFFF;
rommem[22164] <= 16'hFFFF;
rommem[22165] <= 16'hFFFF;
rommem[22166] <= 16'hFFFF;
rommem[22167] <= 16'hFFFF;
rommem[22168] <= 16'hFFFF;
rommem[22169] <= 16'hFFFF;
rommem[22170] <= 16'hFFFF;
rommem[22171] <= 16'hFFFF;
rommem[22172] <= 16'hFFFF;
rommem[22173] <= 16'hFFFF;
rommem[22174] <= 16'hFFFF;
rommem[22175] <= 16'hFFFF;
rommem[22176] <= 16'hFFFF;
rommem[22177] <= 16'hFFFF;
rommem[22178] <= 16'hFFFF;
rommem[22179] <= 16'hFFFF;
rommem[22180] <= 16'hFFFF;
rommem[22181] <= 16'hFFFF;
rommem[22182] <= 16'hFFFF;
rommem[22183] <= 16'hFFFF;
rommem[22184] <= 16'hFFFF;
rommem[22185] <= 16'hFFFF;
rommem[22186] <= 16'hFFFF;
rommem[22187] <= 16'hFFFF;
rommem[22188] <= 16'hFFFF;
rommem[22189] <= 16'hFFFF;
rommem[22190] <= 16'hFFFF;
rommem[22191] <= 16'hFFFF;
rommem[22192] <= 16'hFFFF;
rommem[22193] <= 16'hFFFF;
rommem[22194] <= 16'hFFFF;
rommem[22195] <= 16'hFFFF;
rommem[22196] <= 16'hFFFF;
rommem[22197] <= 16'hFFFF;
rommem[22198] <= 16'hFFFF;
rommem[22199] <= 16'hFFFF;
rommem[22200] <= 16'hFFFF;
rommem[22201] <= 16'hFFFF;
rommem[22202] <= 16'hFFFF;
rommem[22203] <= 16'hFFFF;
rommem[22204] <= 16'hFFFF;
rommem[22205] <= 16'hFFFF;
rommem[22206] <= 16'hFFFF;
rommem[22207] <= 16'hFFFF;
rommem[22208] <= 16'hFFFF;
rommem[22209] <= 16'hFFFF;
rommem[22210] <= 16'hFFFF;
rommem[22211] <= 16'hFFFF;
rommem[22212] <= 16'hFFFF;
rommem[22213] <= 16'hFFFF;
rommem[22214] <= 16'hFFFF;
rommem[22215] <= 16'hFFFF;
rommem[22216] <= 16'hFFFF;
rommem[22217] <= 16'hFFFF;
rommem[22218] <= 16'hFFFF;
rommem[22219] <= 16'hFFFF;
rommem[22220] <= 16'hFFFF;
rommem[22221] <= 16'hFFFF;
rommem[22222] <= 16'hFFFF;
rommem[22223] <= 16'hFFFF;
rommem[22224] <= 16'hFFFF;
rommem[22225] <= 16'hFFFF;
rommem[22226] <= 16'hFFFF;
rommem[22227] <= 16'hFFFF;
rommem[22228] <= 16'hFFFF;
rommem[22229] <= 16'hFFFF;
rommem[22230] <= 16'hFFFF;
rommem[22231] <= 16'hFFFF;
rommem[22232] <= 16'hFFFF;
rommem[22233] <= 16'hFFFF;
rommem[22234] <= 16'hFFFF;
rommem[22235] <= 16'hFFFF;
rommem[22236] <= 16'hFFFF;
rommem[22237] <= 16'hFFFF;
rommem[22238] <= 16'hFFFF;
rommem[22239] <= 16'hFFFF;
rommem[22240] <= 16'hFFFF;
rommem[22241] <= 16'hFFFF;
rommem[22242] <= 16'hFFFF;
rommem[22243] <= 16'hFFFF;
rommem[22244] <= 16'hFFFF;
rommem[22245] <= 16'hFFFF;
rommem[22246] <= 16'hFFFF;
rommem[22247] <= 16'hFFFF;
rommem[22248] <= 16'hFFFF;
rommem[22249] <= 16'hFFFF;
rommem[22250] <= 16'hFFFF;
rommem[22251] <= 16'hFFFF;
rommem[22252] <= 16'hFFFF;
rommem[22253] <= 16'hFFFF;
rommem[22254] <= 16'hFFFF;
rommem[22255] <= 16'hFFFF;
rommem[22256] <= 16'hFFFF;
rommem[22257] <= 16'hFFFF;
rommem[22258] <= 16'hFFFF;
rommem[22259] <= 16'hFFFF;
rommem[22260] <= 16'hFFFF;
rommem[22261] <= 16'hFFFF;
rommem[22262] <= 16'hFFFF;
rommem[22263] <= 16'hFFFF;
rommem[22264] <= 16'hFFFF;
rommem[22265] <= 16'hFFFF;
rommem[22266] <= 16'hFFFF;
rommem[22267] <= 16'hFFFF;
rommem[22268] <= 16'hFFFF;
rommem[22269] <= 16'hFFFF;
rommem[22270] <= 16'hFFFF;
rommem[22271] <= 16'hFFFF;
rommem[22272] <= 16'hFFFF;
rommem[22273] <= 16'hFFFF;
rommem[22274] <= 16'hFFFF;
rommem[22275] <= 16'hFFFF;
rommem[22276] <= 16'hFFFF;
rommem[22277] <= 16'hFFFF;
rommem[22278] <= 16'hFFFF;
rommem[22279] <= 16'hFFFF;
rommem[22280] <= 16'hFFFF;
rommem[22281] <= 16'hFFFF;
rommem[22282] <= 16'hFFFF;
rommem[22283] <= 16'hFFFF;
rommem[22284] <= 16'hFFFF;
rommem[22285] <= 16'hFFFF;
rommem[22286] <= 16'hFFFF;
rommem[22287] <= 16'hFFFF;
rommem[22288] <= 16'hFFFF;
rommem[22289] <= 16'hFFFF;
rommem[22290] <= 16'hFFFF;
rommem[22291] <= 16'hFFFF;
rommem[22292] <= 16'hFFFF;
rommem[22293] <= 16'hFFFF;
rommem[22294] <= 16'hFFFF;
rommem[22295] <= 16'hFFFF;
rommem[22296] <= 16'hFFFF;
rommem[22297] <= 16'hFFFF;
rommem[22298] <= 16'hFFFF;
rommem[22299] <= 16'hFFFF;
rommem[22300] <= 16'hFFFF;
rommem[22301] <= 16'hFFFF;
rommem[22302] <= 16'hFFFF;
rommem[22303] <= 16'hFFFF;
rommem[22304] <= 16'hFFFF;
rommem[22305] <= 16'hFFFF;
rommem[22306] <= 16'hFFFF;
rommem[22307] <= 16'hFFFF;
rommem[22308] <= 16'hFFFF;
rommem[22309] <= 16'hFFFF;
rommem[22310] <= 16'hFFFF;
rommem[22311] <= 16'hFFFF;
rommem[22312] <= 16'hFFFF;
rommem[22313] <= 16'hFFFF;
rommem[22314] <= 16'hFFFF;
rommem[22315] <= 16'hFFFF;
rommem[22316] <= 16'hFFFF;
rommem[22317] <= 16'hFFFF;
rommem[22318] <= 16'hFFFF;
rommem[22319] <= 16'hFFFF;
rommem[22320] <= 16'hFFFF;
rommem[22321] <= 16'hFFFF;
rommem[22322] <= 16'hFFFF;
rommem[22323] <= 16'hFFFF;
rommem[22324] <= 16'hFFFF;
rommem[22325] <= 16'hFFFF;
rommem[22326] <= 16'hFFFF;
rommem[22327] <= 16'hFFFF;
rommem[22328] <= 16'hFFFF;
rommem[22329] <= 16'hFFFF;
rommem[22330] <= 16'hFFFF;
rommem[22331] <= 16'hFFFF;
rommem[22332] <= 16'hFFFF;
rommem[22333] <= 16'hFFFF;
rommem[22334] <= 16'hFFFF;
rommem[22335] <= 16'hFFFF;
rommem[22336] <= 16'hFFFF;
rommem[22337] <= 16'hFFFF;
rommem[22338] <= 16'hFFFF;
rommem[22339] <= 16'hFFFF;
rommem[22340] <= 16'hFFFF;
rommem[22341] <= 16'hFFFF;
rommem[22342] <= 16'hFFFF;
rommem[22343] <= 16'hFFFF;
rommem[22344] <= 16'hFFFF;
rommem[22345] <= 16'hFFFF;
rommem[22346] <= 16'hFFFF;
rommem[22347] <= 16'hFFFF;
rommem[22348] <= 16'hFFFF;
rommem[22349] <= 16'hFFFF;
rommem[22350] <= 16'hFFFF;
rommem[22351] <= 16'hFFFF;
rommem[22352] <= 16'hFFFF;
rommem[22353] <= 16'hFFFF;
rommem[22354] <= 16'hFFFF;
rommem[22355] <= 16'hFFFF;
rommem[22356] <= 16'hFFFF;
rommem[22357] <= 16'hFFFF;
rommem[22358] <= 16'hFFFF;
rommem[22359] <= 16'hFFFF;
rommem[22360] <= 16'hFFFF;
rommem[22361] <= 16'hFFFF;
rommem[22362] <= 16'hFFFF;
rommem[22363] <= 16'hFFFF;
rommem[22364] <= 16'hFFFF;
rommem[22365] <= 16'hFFFF;
rommem[22366] <= 16'hFFFF;
rommem[22367] <= 16'hFFFF;
rommem[22368] <= 16'hFFFF;
rommem[22369] <= 16'hFFFF;
rommem[22370] <= 16'hFFFF;
rommem[22371] <= 16'hFFFF;
rommem[22372] <= 16'hFFFF;
rommem[22373] <= 16'hFFFF;
rommem[22374] <= 16'hFFFF;
rommem[22375] <= 16'hFFFF;
rommem[22376] <= 16'hFFFF;
rommem[22377] <= 16'hFFFF;
rommem[22378] <= 16'hFFFF;
rommem[22379] <= 16'hFFFF;
rommem[22380] <= 16'hFFFF;
rommem[22381] <= 16'hFFFF;
rommem[22382] <= 16'hFFFF;
rommem[22383] <= 16'hFFFF;
rommem[22384] <= 16'hFFFF;
rommem[22385] <= 16'hFFFF;
rommem[22386] <= 16'hFFFF;
rommem[22387] <= 16'hFFFF;
rommem[22388] <= 16'hFFFF;
rommem[22389] <= 16'hFFFF;
rommem[22390] <= 16'hFFFF;
rommem[22391] <= 16'hFFFF;
rommem[22392] <= 16'hFFFF;
rommem[22393] <= 16'hFFFF;
rommem[22394] <= 16'hFFFF;
rommem[22395] <= 16'hFFFF;
rommem[22396] <= 16'hFFFF;
rommem[22397] <= 16'hFFFF;
rommem[22398] <= 16'hFFFF;
rommem[22399] <= 16'hFFFF;
rommem[22400] <= 16'hFFFF;
rommem[22401] <= 16'hFFFF;
rommem[22402] <= 16'hFFFF;
rommem[22403] <= 16'hFFFF;
rommem[22404] <= 16'hFFFF;
rommem[22405] <= 16'hFFFF;
rommem[22406] <= 16'hFFFF;
rommem[22407] <= 16'hFFFF;
rommem[22408] <= 16'hFFFF;
rommem[22409] <= 16'hFFFF;
rommem[22410] <= 16'hFFFF;
rommem[22411] <= 16'hFFFF;
rommem[22412] <= 16'hFFFF;
rommem[22413] <= 16'hFFFF;
rommem[22414] <= 16'hFFFF;
rommem[22415] <= 16'hFFFF;
rommem[22416] <= 16'hFFFF;
rommem[22417] <= 16'hFFFF;
rommem[22418] <= 16'hFFFF;
rommem[22419] <= 16'hFFFF;
rommem[22420] <= 16'hFFFF;
rommem[22421] <= 16'hFFFF;
rommem[22422] <= 16'hFFFF;
rommem[22423] <= 16'hFFFF;
rommem[22424] <= 16'hFFFF;
rommem[22425] <= 16'hFFFF;
rommem[22426] <= 16'hFFFF;
rommem[22427] <= 16'hFFFF;
rommem[22428] <= 16'hFFFF;
rommem[22429] <= 16'hFFFF;
rommem[22430] <= 16'hFFFF;
rommem[22431] <= 16'hFFFF;
rommem[22432] <= 16'hFFFF;
rommem[22433] <= 16'hFFFF;
rommem[22434] <= 16'hFFFF;
rommem[22435] <= 16'hFFFF;
rommem[22436] <= 16'hFFFF;
rommem[22437] <= 16'hFFFF;
rommem[22438] <= 16'hFFFF;
rommem[22439] <= 16'hFFFF;
rommem[22440] <= 16'hFFFF;
rommem[22441] <= 16'hFFFF;
rommem[22442] <= 16'hFFFF;
rommem[22443] <= 16'hFFFF;
rommem[22444] <= 16'hFFFF;
rommem[22445] <= 16'hFFFF;
rommem[22446] <= 16'hFFFF;
rommem[22447] <= 16'hFFFF;
rommem[22448] <= 16'hFFFF;
rommem[22449] <= 16'hFFFF;
rommem[22450] <= 16'hFFFF;
rommem[22451] <= 16'hFFFF;
rommem[22452] <= 16'hFFFF;
rommem[22453] <= 16'hFFFF;
rommem[22454] <= 16'hFFFF;
rommem[22455] <= 16'hFFFF;
rommem[22456] <= 16'hFFFF;
rommem[22457] <= 16'hFFFF;
rommem[22458] <= 16'hFFFF;
rommem[22459] <= 16'hFFFF;
rommem[22460] <= 16'hFFFF;
rommem[22461] <= 16'hFFFF;
rommem[22462] <= 16'hFFFF;
rommem[22463] <= 16'hFFFF;
rommem[22464] <= 16'hFFFF;
rommem[22465] <= 16'hFFFF;
rommem[22466] <= 16'hFFFF;
rommem[22467] <= 16'hFFFF;
rommem[22468] <= 16'hFFFF;
rommem[22469] <= 16'hFFFF;
rommem[22470] <= 16'hFFFF;
rommem[22471] <= 16'hFFFF;
rommem[22472] <= 16'hFFFF;
rommem[22473] <= 16'hFFFF;
rommem[22474] <= 16'hFFFF;
rommem[22475] <= 16'hFFFF;
rommem[22476] <= 16'hFFFF;
rommem[22477] <= 16'hFFFF;
rommem[22478] <= 16'hFFFF;
rommem[22479] <= 16'hFFFF;
rommem[22480] <= 16'hFFFF;
rommem[22481] <= 16'hFFFF;
rommem[22482] <= 16'hFFFF;
rommem[22483] <= 16'hFFFF;
rommem[22484] <= 16'hFFFF;
rommem[22485] <= 16'hFFFF;
rommem[22486] <= 16'hFFFF;
rommem[22487] <= 16'hFFFF;
rommem[22488] <= 16'hFFFF;
rommem[22489] <= 16'hFFFF;
rommem[22490] <= 16'hFFFF;
rommem[22491] <= 16'hFFFF;
rommem[22492] <= 16'hFFFF;
rommem[22493] <= 16'hFFFF;
rommem[22494] <= 16'hFFFF;
rommem[22495] <= 16'hFFFF;
rommem[22496] <= 16'hFFFF;
rommem[22497] <= 16'hFFFF;
rommem[22498] <= 16'hFFFF;
rommem[22499] <= 16'hFFFF;
rommem[22500] <= 16'hFFFF;
rommem[22501] <= 16'hFFFF;
rommem[22502] <= 16'hFFFF;
rommem[22503] <= 16'hFFFF;
rommem[22504] <= 16'hFFFF;
rommem[22505] <= 16'hFFFF;
rommem[22506] <= 16'hFFFF;
rommem[22507] <= 16'hFFFF;
rommem[22508] <= 16'hFFFF;
rommem[22509] <= 16'hFFFF;
rommem[22510] <= 16'hFFFF;
rommem[22511] <= 16'hFFFF;
rommem[22512] <= 16'hFFFF;
rommem[22513] <= 16'hFFFF;
rommem[22514] <= 16'hFFFF;
rommem[22515] <= 16'hFFFF;
rommem[22516] <= 16'hFFFF;
rommem[22517] <= 16'hFFFF;
rommem[22518] <= 16'hFFFF;
rommem[22519] <= 16'hFFFF;
rommem[22520] <= 16'hFFFF;
rommem[22521] <= 16'hFFFF;
rommem[22522] <= 16'hFFFF;
rommem[22523] <= 16'hFFFF;
rommem[22524] <= 16'hFFFF;
rommem[22525] <= 16'hFFFF;
rommem[22526] <= 16'hFFFF;
rommem[22527] <= 16'hFFFF;
rommem[22528] <= 16'hFFFF;
rommem[22529] <= 16'hFFFF;
rommem[22530] <= 16'hFFFF;
rommem[22531] <= 16'hFFFF;
rommem[22532] <= 16'hFFFF;
rommem[22533] <= 16'hFFFF;
rommem[22534] <= 16'hFFFF;
rommem[22535] <= 16'hFFFF;
rommem[22536] <= 16'hFFFF;
rommem[22537] <= 16'hFFFF;
rommem[22538] <= 16'hFFFF;
rommem[22539] <= 16'hFFFF;
rommem[22540] <= 16'hFFFF;
rommem[22541] <= 16'hFFFF;
rommem[22542] <= 16'hFFFF;
rommem[22543] <= 16'hFFFF;
rommem[22544] <= 16'hFFFF;
rommem[22545] <= 16'hFFFF;
rommem[22546] <= 16'hFFFF;
rommem[22547] <= 16'hFFFF;
rommem[22548] <= 16'hFFFF;
rommem[22549] <= 16'hFFFF;
rommem[22550] <= 16'hFFFF;
rommem[22551] <= 16'hFFFF;
rommem[22552] <= 16'hFFFF;
rommem[22553] <= 16'hFFFF;
rommem[22554] <= 16'hFFFF;
rommem[22555] <= 16'hFFFF;
rommem[22556] <= 16'hFFFF;
rommem[22557] <= 16'hFFFF;
rommem[22558] <= 16'hFFFF;
rommem[22559] <= 16'hFFFF;
rommem[22560] <= 16'hFFFF;
rommem[22561] <= 16'hFFFF;
rommem[22562] <= 16'hFFFF;
rommem[22563] <= 16'hFFFF;
rommem[22564] <= 16'hFFFF;
rommem[22565] <= 16'hFFFF;
rommem[22566] <= 16'hFFFF;
rommem[22567] <= 16'hFFFF;
rommem[22568] <= 16'hFFFF;
rommem[22569] <= 16'hFFFF;
rommem[22570] <= 16'hFFFF;
rommem[22571] <= 16'hFFFF;
rommem[22572] <= 16'hFFFF;
rommem[22573] <= 16'hFFFF;
rommem[22574] <= 16'hFFFF;
rommem[22575] <= 16'hFFFF;
rommem[22576] <= 16'hFFFF;
rommem[22577] <= 16'hFFFF;
rommem[22578] <= 16'hFFFF;
rommem[22579] <= 16'hFFFF;
rommem[22580] <= 16'hFFFF;
rommem[22581] <= 16'hFFFF;
rommem[22582] <= 16'hFFFF;
rommem[22583] <= 16'hFFFF;
rommem[22584] <= 16'hFFFF;
rommem[22585] <= 16'hFFFF;
rommem[22586] <= 16'hFFFF;
rommem[22587] <= 16'hFFFF;
rommem[22588] <= 16'hFFFF;
rommem[22589] <= 16'hFFFF;
rommem[22590] <= 16'hFFFF;
rommem[22591] <= 16'hFFFF;
rommem[22592] <= 16'hFFFF;
rommem[22593] <= 16'hFFFF;
rommem[22594] <= 16'hFFFF;
rommem[22595] <= 16'hFFFF;
rommem[22596] <= 16'hFFFF;
rommem[22597] <= 16'hFFFF;
rommem[22598] <= 16'hFFFF;
rommem[22599] <= 16'hFFFF;
rommem[22600] <= 16'hFFFF;
rommem[22601] <= 16'hFFFF;
rommem[22602] <= 16'hFFFF;
rommem[22603] <= 16'hFFFF;
rommem[22604] <= 16'hFFFF;
rommem[22605] <= 16'hFFFF;
rommem[22606] <= 16'hFFFF;
rommem[22607] <= 16'hFFFF;
rommem[22608] <= 16'hFFFF;
rommem[22609] <= 16'hFFFF;
rommem[22610] <= 16'hFFFF;
rommem[22611] <= 16'hFFFF;
rommem[22612] <= 16'hFFFF;
rommem[22613] <= 16'hFFFF;
rommem[22614] <= 16'hFFFF;
rommem[22615] <= 16'hFFFF;
rommem[22616] <= 16'hFFFF;
rommem[22617] <= 16'hFFFF;
rommem[22618] <= 16'hFFFF;
rommem[22619] <= 16'hFFFF;
rommem[22620] <= 16'hFFFF;
rommem[22621] <= 16'hFFFF;
rommem[22622] <= 16'hFFFF;
rommem[22623] <= 16'hFFFF;
rommem[22624] <= 16'hFFFF;
rommem[22625] <= 16'hFFFF;
rommem[22626] <= 16'hFFFF;
rommem[22627] <= 16'hFFFF;
rommem[22628] <= 16'hFFFF;
rommem[22629] <= 16'hFFFF;
rommem[22630] <= 16'hFFFF;
rommem[22631] <= 16'hFFFF;
rommem[22632] <= 16'hFFFF;
rommem[22633] <= 16'hFFFF;
rommem[22634] <= 16'hFFFF;
rommem[22635] <= 16'hFFFF;
rommem[22636] <= 16'hFFFF;
rommem[22637] <= 16'hFFFF;
rommem[22638] <= 16'hFFFF;
rommem[22639] <= 16'hFFFF;
rommem[22640] <= 16'hFFFF;
rommem[22641] <= 16'hFFFF;
rommem[22642] <= 16'hFFFF;
rommem[22643] <= 16'hFFFF;
rommem[22644] <= 16'hFFFF;
rommem[22645] <= 16'hFFFF;
rommem[22646] <= 16'hFFFF;
rommem[22647] <= 16'hFFFF;
rommem[22648] <= 16'hFFFF;
rommem[22649] <= 16'hFFFF;
rommem[22650] <= 16'hFFFF;
rommem[22651] <= 16'hFFFF;
rommem[22652] <= 16'hFFFF;
rommem[22653] <= 16'hFFFF;
rommem[22654] <= 16'hFFFF;
rommem[22655] <= 16'hFFFF;
rommem[22656] <= 16'hFFFF;
rommem[22657] <= 16'hFFFF;
rommem[22658] <= 16'hFFFF;
rommem[22659] <= 16'hFFFF;
rommem[22660] <= 16'hFFFF;
rommem[22661] <= 16'hFFFF;
rommem[22662] <= 16'hFFFF;
rommem[22663] <= 16'hFFFF;
rommem[22664] <= 16'hFFFF;
rommem[22665] <= 16'hFFFF;
rommem[22666] <= 16'hFFFF;
rommem[22667] <= 16'hFFFF;
rommem[22668] <= 16'hFFFF;
rommem[22669] <= 16'hFFFF;
rommem[22670] <= 16'hFFFF;
rommem[22671] <= 16'hFFFF;
rommem[22672] <= 16'hFFFF;
rommem[22673] <= 16'hFFFF;
rommem[22674] <= 16'hFFFF;
rommem[22675] <= 16'hFFFF;
rommem[22676] <= 16'hFFFF;
rommem[22677] <= 16'hFFFF;
rommem[22678] <= 16'hFFFF;
rommem[22679] <= 16'hFFFF;
rommem[22680] <= 16'hFFFF;
rommem[22681] <= 16'hFFFF;
rommem[22682] <= 16'hFFFF;
rommem[22683] <= 16'hFFFF;
rommem[22684] <= 16'hFFFF;
rommem[22685] <= 16'hFFFF;
rommem[22686] <= 16'hFFFF;
rommem[22687] <= 16'hFFFF;
rommem[22688] <= 16'hFFFF;
rommem[22689] <= 16'hFFFF;
rommem[22690] <= 16'hFFFF;
rommem[22691] <= 16'hFFFF;
rommem[22692] <= 16'hFFFF;
rommem[22693] <= 16'hFFFF;
rommem[22694] <= 16'hFFFF;
rommem[22695] <= 16'hFFFF;
rommem[22696] <= 16'hFFFF;
rommem[22697] <= 16'hFFFF;
rommem[22698] <= 16'hFFFF;
rommem[22699] <= 16'hFFFF;
rommem[22700] <= 16'hFFFF;
rommem[22701] <= 16'hFFFF;
rommem[22702] <= 16'hFFFF;
rommem[22703] <= 16'hFFFF;
rommem[22704] <= 16'hFFFF;
rommem[22705] <= 16'hFFFF;
rommem[22706] <= 16'hFFFF;
rommem[22707] <= 16'hFFFF;
rommem[22708] <= 16'hFFFF;
rommem[22709] <= 16'hFFFF;
rommem[22710] <= 16'hFFFF;
rommem[22711] <= 16'hFFFF;
rommem[22712] <= 16'hFFFF;
rommem[22713] <= 16'hFFFF;
rommem[22714] <= 16'hFFFF;
rommem[22715] <= 16'hFFFF;
rommem[22716] <= 16'hFFFF;
rommem[22717] <= 16'hFFFF;
rommem[22718] <= 16'hFFFF;
rommem[22719] <= 16'hFFFF;
rommem[22720] <= 16'hFFFF;
rommem[22721] <= 16'hFFFF;
rommem[22722] <= 16'hFFFF;
rommem[22723] <= 16'hFFFF;
rommem[22724] <= 16'hFFFF;
rommem[22725] <= 16'hFFFF;
rommem[22726] <= 16'hFFFF;
rommem[22727] <= 16'hFFFF;
rommem[22728] <= 16'hFFFF;
rommem[22729] <= 16'hFFFF;
rommem[22730] <= 16'hFFFF;
rommem[22731] <= 16'hFFFF;
rommem[22732] <= 16'hFFFF;
rommem[22733] <= 16'hFFFF;
rommem[22734] <= 16'hFFFF;
rommem[22735] <= 16'hFFFF;
rommem[22736] <= 16'hFFFF;
rommem[22737] <= 16'hFFFF;
rommem[22738] <= 16'hFFFF;
rommem[22739] <= 16'hFFFF;
rommem[22740] <= 16'hFFFF;
rommem[22741] <= 16'hFFFF;
rommem[22742] <= 16'hFFFF;
rommem[22743] <= 16'hFFFF;
rommem[22744] <= 16'hFFFF;
rommem[22745] <= 16'hFFFF;
rommem[22746] <= 16'hFFFF;
rommem[22747] <= 16'hFFFF;
rommem[22748] <= 16'hFFFF;
rommem[22749] <= 16'hFFFF;
rommem[22750] <= 16'hFFFF;
rommem[22751] <= 16'hFFFF;
rommem[22752] <= 16'hFFFF;
rommem[22753] <= 16'hFFFF;
rommem[22754] <= 16'hFFFF;
rommem[22755] <= 16'hFFFF;
rommem[22756] <= 16'hFFFF;
rommem[22757] <= 16'hFFFF;
rommem[22758] <= 16'hFFFF;
rommem[22759] <= 16'hFFFF;
rommem[22760] <= 16'hFFFF;
rommem[22761] <= 16'hFFFF;
rommem[22762] <= 16'hFFFF;
rommem[22763] <= 16'hFFFF;
rommem[22764] <= 16'hFFFF;
rommem[22765] <= 16'hFFFF;
rommem[22766] <= 16'hFFFF;
rommem[22767] <= 16'hFFFF;
rommem[22768] <= 16'hFFFF;
rommem[22769] <= 16'hFFFF;
rommem[22770] <= 16'hFFFF;
rommem[22771] <= 16'hFFFF;
rommem[22772] <= 16'hFFFF;
rommem[22773] <= 16'hFFFF;
rommem[22774] <= 16'hFFFF;
rommem[22775] <= 16'hFFFF;
rommem[22776] <= 16'hFFFF;
rommem[22777] <= 16'hFFFF;
rommem[22778] <= 16'hFFFF;
rommem[22779] <= 16'hFFFF;
rommem[22780] <= 16'hFFFF;
rommem[22781] <= 16'hFFFF;
rommem[22782] <= 16'hFFFF;
rommem[22783] <= 16'hFFFF;
rommem[22784] <= 16'hFFFF;
rommem[22785] <= 16'hFFFF;
rommem[22786] <= 16'hFFFF;
rommem[22787] <= 16'hFFFF;
rommem[22788] <= 16'hFFFF;
rommem[22789] <= 16'hFFFF;
rommem[22790] <= 16'hFFFF;
rommem[22791] <= 16'hFFFF;
rommem[22792] <= 16'hFFFF;
rommem[22793] <= 16'hFFFF;
rommem[22794] <= 16'hFFFF;
rommem[22795] <= 16'hFFFF;
rommem[22796] <= 16'hFFFF;
rommem[22797] <= 16'hFFFF;
rommem[22798] <= 16'hFFFF;
rommem[22799] <= 16'hFFFF;
rommem[22800] <= 16'hFFFF;
rommem[22801] <= 16'hFFFF;
rommem[22802] <= 16'hFFFF;
rommem[22803] <= 16'hFFFF;
rommem[22804] <= 16'hFFFF;
rommem[22805] <= 16'hFFFF;
rommem[22806] <= 16'hFFFF;
rommem[22807] <= 16'hFFFF;
rommem[22808] <= 16'hFFFF;
rommem[22809] <= 16'hFFFF;
rommem[22810] <= 16'hFFFF;
rommem[22811] <= 16'hFFFF;
rommem[22812] <= 16'hFFFF;
rommem[22813] <= 16'hFFFF;
rommem[22814] <= 16'hFFFF;
rommem[22815] <= 16'hFFFF;
rommem[22816] <= 16'hFFFF;
rommem[22817] <= 16'hFFFF;
rommem[22818] <= 16'hFFFF;
rommem[22819] <= 16'hFFFF;
rommem[22820] <= 16'hFFFF;
rommem[22821] <= 16'hFFFF;
rommem[22822] <= 16'hFFFF;
rommem[22823] <= 16'hFFFF;
rommem[22824] <= 16'hFFFF;
rommem[22825] <= 16'hFFFF;
rommem[22826] <= 16'hFFFF;
rommem[22827] <= 16'hFFFF;
rommem[22828] <= 16'hFFFF;
rommem[22829] <= 16'hFFFF;
rommem[22830] <= 16'hFFFF;
rommem[22831] <= 16'hFFFF;
rommem[22832] <= 16'hFFFF;
rommem[22833] <= 16'hFFFF;
rommem[22834] <= 16'hFFFF;
rommem[22835] <= 16'hFFFF;
rommem[22836] <= 16'hFFFF;
rommem[22837] <= 16'hFFFF;
rommem[22838] <= 16'hFFFF;
rommem[22839] <= 16'hFFFF;
rommem[22840] <= 16'hFFFF;
rommem[22841] <= 16'hFFFF;
rommem[22842] <= 16'hFFFF;
rommem[22843] <= 16'hFFFF;
rommem[22844] <= 16'hFFFF;
rommem[22845] <= 16'hFFFF;
rommem[22846] <= 16'hFFFF;
rommem[22847] <= 16'hFFFF;
rommem[22848] <= 16'hFFFF;
rommem[22849] <= 16'hFFFF;
rommem[22850] <= 16'hFFFF;
rommem[22851] <= 16'hFFFF;
rommem[22852] <= 16'hFFFF;
rommem[22853] <= 16'hFFFF;
rommem[22854] <= 16'hFFFF;
rommem[22855] <= 16'hFFFF;
rommem[22856] <= 16'hFFFF;
rommem[22857] <= 16'hFFFF;
rommem[22858] <= 16'hFFFF;
rommem[22859] <= 16'hFFFF;
rommem[22860] <= 16'hFFFF;
rommem[22861] <= 16'hFFFF;
rommem[22862] <= 16'hFFFF;
rommem[22863] <= 16'hFFFF;
rommem[22864] <= 16'hFFFF;
rommem[22865] <= 16'hFFFF;
rommem[22866] <= 16'hFFFF;
rommem[22867] <= 16'hFFFF;
rommem[22868] <= 16'hFFFF;
rommem[22869] <= 16'hFFFF;
rommem[22870] <= 16'hFFFF;
rommem[22871] <= 16'hFFFF;
rommem[22872] <= 16'hFFFF;
rommem[22873] <= 16'hFFFF;
rommem[22874] <= 16'hFFFF;
rommem[22875] <= 16'hFFFF;
rommem[22876] <= 16'hFFFF;
rommem[22877] <= 16'hFFFF;
rommem[22878] <= 16'hFFFF;
rommem[22879] <= 16'hFFFF;
rommem[22880] <= 16'hFFFF;
rommem[22881] <= 16'hFFFF;
rommem[22882] <= 16'hFFFF;
rommem[22883] <= 16'hFFFF;
rommem[22884] <= 16'hFFFF;
rommem[22885] <= 16'hFFFF;
rommem[22886] <= 16'hFFFF;
rommem[22887] <= 16'hFFFF;
rommem[22888] <= 16'hFFFF;
rommem[22889] <= 16'hFFFF;
rommem[22890] <= 16'hFFFF;
rommem[22891] <= 16'hFFFF;
rommem[22892] <= 16'hFFFF;
rommem[22893] <= 16'hFFFF;
rommem[22894] <= 16'hFFFF;
rommem[22895] <= 16'hFFFF;
rommem[22896] <= 16'hFFFF;
rommem[22897] <= 16'hFFFF;
rommem[22898] <= 16'hFFFF;
rommem[22899] <= 16'hFFFF;
rommem[22900] <= 16'hFFFF;
rommem[22901] <= 16'hFFFF;
rommem[22902] <= 16'hFFFF;
rommem[22903] <= 16'hFFFF;
rommem[22904] <= 16'hFFFF;
rommem[22905] <= 16'hFFFF;
rommem[22906] <= 16'hFFFF;
rommem[22907] <= 16'hFFFF;
rommem[22908] <= 16'hFFFF;
rommem[22909] <= 16'hFFFF;
rommem[22910] <= 16'hFFFF;
rommem[22911] <= 16'hFFFF;
rommem[22912] <= 16'hFFFF;
rommem[22913] <= 16'hFFFF;
rommem[22914] <= 16'hFFFF;
rommem[22915] <= 16'hFFFF;
rommem[22916] <= 16'hFFFF;
rommem[22917] <= 16'hFFFF;
rommem[22918] <= 16'hFFFF;
rommem[22919] <= 16'hFFFF;
rommem[22920] <= 16'hFFFF;
rommem[22921] <= 16'hFFFF;
rommem[22922] <= 16'hFFFF;
rommem[22923] <= 16'hFFFF;
rommem[22924] <= 16'hFFFF;
rommem[22925] <= 16'hFFFF;
rommem[22926] <= 16'hFFFF;
rommem[22927] <= 16'hFFFF;
rommem[22928] <= 16'hFFFF;
rommem[22929] <= 16'hFFFF;
rommem[22930] <= 16'hFFFF;
rommem[22931] <= 16'hFFFF;
rommem[22932] <= 16'hFFFF;
rommem[22933] <= 16'hFFFF;
rommem[22934] <= 16'hFFFF;
rommem[22935] <= 16'hFFFF;
rommem[22936] <= 16'hFFFF;
rommem[22937] <= 16'hFFFF;
rommem[22938] <= 16'hFFFF;
rommem[22939] <= 16'hFFFF;
rommem[22940] <= 16'hFFFF;
rommem[22941] <= 16'hFFFF;
rommem[22942] <= 16'hFFFF;
rommem[22943] <= 16'hFFFF;
rommem[22944] <= 16'hFFFF;
rommem[22945] <= 16'hFFFF;
rommem[22946] <= 16'hFFFF;
rommem[22947] <= 16'hFFFF;
rommem[22948] <= 16'hFFFF;
rommem[22949] <= 16'hFFFF;
rommem[22950] <= 16'hFFFF;
rommem[22951] <= 16'hFFFF;
rommem[22952] <= 16'hFFFF;
rommem[22953] <= 16'hFFFF;
rommem[22954] <= 16'hFFFF;
rommem[22955] <= 16'hFFFF;
rommem[22956] <= 16'hFFFF;
rommem[22957] <= 16'hFFFF;
rommem[22958] <= 16'hFFFF;
rommem[22959] <= 16'hFFFF;
rommem[22960] <= 16'hFFFF;
rommem[22961] <= 16'hFFFF;
rommem[22962] <= 16'hFFFF;
rommem[22963] <= 16'hFFFF;
rommem[22964] <= 16'hFFFF;
rommem[22965] <= 16'hFFFF;
rommem[22966] <= 16'hFFFF;
rommem[22967] <= 16'hFFFF;
rommem[22968] <= 16'hFFFF;
rommem[22969] <= 16'hFFFF;
rommem[22970] <= 16'hFFFF;
rommem[22971] <= 16'hFFFF;
rommem[22972] <= 16'hFFFF;
rommem[22973] <= 16'hFFFF;
rommem[22974] <= 16'hFFFF;
rommem[22975] <= 16'hFFFF;
rommem[22976] <= 16'hFFFF;
rommem[22977] <= 16'hFFFF;
rommem[22978] <= 16'hFFFF;
rommem[22979] <= 16'hFFFF;
rommem[22980] <= 16'hFFFF;
rommem[22981] <= 16'hFFFF;
rommem[22982] <= 16'hFFFF;
rommem[22983] <= 16'hFFFF;
rommem[22984] <= 16'hFFFF;
rommem[22985] <= 16'hFFFF;
rommem[22986] <= 16'hFFFF;
rommem[22987] <= 16'hFFFF;
rommem[22988] <= 16'hFFFF;
rommem[22989] <= 16'hFFFF;
rommem[22990] <= 16'hFFFF;
rommem[22991] <= 16'hFFFF;
rommem[22992] <= 16'hFFFF;
rommem[22993] <= 16'hFFFF;
rommem[22994] <= 16'hFFFF;
rommem[22995] <= 16'hFFFF;
rommem[22996] <= 16'hFFFF;
rommem[22997] <= 16'hFFFF;
rommem[22998] <= 16'hFFFF;
rommem[22999] <= 16'hFFFF;
rommem[23000] <= 16'hFFFF;
rommem[23001] <= 16'hFFFF;
rommem[23002] <= 16'hFFFF;
rommem[23003] <= 16'hFFFF;
rommem[23004] <= 16'hFFFF;
rommem[23005] <= 16'hFFFF;
rommem[23006] <= 16'hFFFF;
rommem[23007] <= 16'hFFFF;
rommem[23008] <= 16'hFFFF;
rommem[23009] <= 16'hFFFF;
rommem[23010] <= 16'hFFFF;
rommem[23011] <= 16'hFFFF;
rommem[23012] <= 16'hFFFF;
rommem[23013] <= 16'hFFFF;
rommem[23014] <= 16'hFFFF;
rommem[23015] <= 16'hFFFF;
rommem[23016] <= 16'hFFFF;
rommem[23017] <= 16'hFFFF;
rommem[23018] <= 16'hFFFF;
rommem[23019] <= 16'hFFFF;
rommem[23020] <= 16'hFFFF;
rommem[23021] <= 16'hFFFF;
rommem[23022] <= 16'hFFFF;
rommem[23023] <= 16'hFFFF;
rommem[23024] <= 16'hFFFF;
rommem[23025] <= 16'hFFFF;
rommem[23026] <= 16'hFFFF;
rommem[23027] <= 16'hFFFF;
rommem[23028] <= 16'hFFFF;
rommem[23029] <= 16'hFFFF;
rommem[23030] <= 16'hFFFF;
rommem[23031] <= 16'hFFFF;
rommem[23032] <= 16'hFFFF;
rommem[23033] <= 16'hFFFF;
rommem[23034] <= 16'hFFFF;
rommem[23035] <= 16'hFFFF;
rommem[23036] <= 16'hFFFF;
rommem[23037] <= 16'hFFFF;
rommem[23038] <= 16'hFFFF;
rommem[23039] <= 16'hFFFF;
rommem[23040] <= 16'hFFFF;
rommem[23041] <= 16'hFFFF;
rommem[23042] <= 16'hFFFF;
rommem[23043] <= 16'hFFFF;
rommem[23044] <= 16'hFFFF;
rommem[23045] <= 16'hFFFF;
rommem[23046] <= 16'hFFFF;
rommem[23047] <= 16'hFFFF;
rommem[23048] <= 16'hFFFF;
rommem[23049] <= 16'hFFFF;
rommem[23050] <= 16'hFFFF;
rommem[23051] <= 16'hFFFF;
rommem[23052] <= 16'hFFFF;
rommem[23053] <= 16'hFFFF;
rommem[23054] <= 16'hFFFF;
rommem[23055] <= 16'hFFFF;
rommem[23056] <= 16'hFFFF;
rommem[23057] <= 16'hFFFF;
rommem[23058] <= 16'hFFFF;
rommem[23059] <= 16'hFFFF;
rommem[23060] <= 16'hFFFF;
rommem[23061] <= 16'hFFFF;
rommem[23062] <= 16'hFFFF;
rommem[23063] <= 16'hFFFF;
rommem[23064] <= 16'hFFFF;
rommem[23065] <= 16'hFFFF;
rommem[23066] <= 16'hFFFF;
rommem[23067] <= 16'hFFFF;
rommem[23068] <= 16'hFFFF;
rommem[23069] <= 16'hFFFF;
rommem[23070] <= 16'hFFFF;
rommem[23071] <= 16'hFFFF;
rommem[23072] <= 16'hFFFF;
rommem[23073] <= 16'hFFFF;
rommem[23074] <= 16'hFFFF;
rommem[23075] <= 16'hFFFF;
rommem[23076] <= 16'hFFFF;
rommem[23077] <= 16'hFFFF;
rommem[23078] <= 16'hFFFF;
rommem[23079] <= 16'hFFFF;
rommem[23080] <= 16'hFFFF;
rommem[23081] <= 16'hFFFF;
rommem[23082] <= 16'hFFFF;
rommem[23083] <= 16'hFFFF;
rommem[23084] <= 16'hFFFF;
rommem[23085] <= 16'hFFFF;
rommem[23086] <= 16'hFFFF;
rommem[23087] <= 16'hFFFF;
rommem[23088] <= 16'hFFFF;
rommem[23089] <= 16'hFFFF;
rommem[23090] <= 16'hFFFF;
rommem[23091] <= 16'hFFFF;
rommem[23092] <= 16'hFFFF;
rommem[23093] <= 16'hFFFF;
rommem[23094] <= 16'hFFFF;
rommem[23095] <= 16'hFFFF;
rommem[23096] <= 16'hFFFF;
rommem[23097] <= 16'hFFFF;
rommem[23098] <= 16'hFFFF;
rommem[23099] <= 16'hFFFF;
rommem[23100] <= 16'hFFFF;
rommem[23101] <= 16'hFFFF;
rommem[23102] <= 16'hFFFF;
rommem[23103] <= 16'hFFFF;
rommem[23104] <= 16'hFFFF;
rommem[23105] <= 16'hFFFF;
rommem[23106] <= 16'hFFFF;
rommem[23107] <= 16'hFFFF;
rommem[23108] <= 16'hFFFF;
rommem[23109] <= 16'hFFFF;
rommem[23110] <= 16'hFFFF;
rommem[23111] <= 16'hFFFF;
rommem[23112] <= 16'hFFFF;
rommem[23113] <= 16'hFFFF;
rommem[23114] <= 16'hFFFF;
rommem[23115] <= 16'hFFFF;
rommem[23116] <= 16'hFFFF;
rommem[23117] <= 16'hFFFF;
rommem[23118] <= 16'hFFFF;
rommem[23119] <= 16'hFFFF;
rommem[23120] <= 16'hFFFF;
rommem[23121] <= 16'hFFFF;
rommem[23122] <= 16'hFFFF;
rommem[23123] <= 16'hFFFF;
rommem[23124] <= 16'hFFFF;
rommem[23125] <= 16'hFFFF;
rommem[23126] <= 16'hFFFF;
rommem[23127] <= 16'hFFFF;
rommem[23128] <= 16'hFFFF;
rommem[23129] <= 16'hFFFF;
rommem[23130] <= 16'hFFFF;
rommem[23131] <= 16'hFFFF;
rommem[23132] <= 16'hFFFF;
rommem[23133] <= 16'hFFFF;
rommem[23134] <= 16'hFFFF;
rommem[23135] <= 16'hFFFF;
rommem[23136] <= 16'hFFFF;
rommem[23137] <= 16'hFFFF;
rommem[23138] <= 16'hFFFF;
rommem[23139] <= 16'hFFFF;
rommem[23140] <= 16'hFFFF;
rommem[23141] <= 16'hFFFF;
rommem[23142] <= 16'hFFFF;
rommem[23143] <= 16'hFFFF;
rommem[23144] <= 16'hFFFF;
rommem[23145] <= 16'hFFFF;
rommem[23146] <= 16'hFFFF;
rommem[23147] <= 16'hFFFF;
rommem[23148] <= 16'hFFFF;
rommem[23149] <= 16'hFFFF;
rommem[23150] <= 16'hFFFF;
rommem[23151] <= 16'hFFFF;
rommem[23152] <= 16'hFFFF;
rommem[23153] <= 16'hFFFF;
rommem[23154] <= 16'hFFFF;
rommem[23155] <= 16'hFFFF;
rommem[23156] <= 16'hFFFF;
rommem[23157] <= 16'hFFFF;
rommem[23158] <= 16'hFFFF;
rommem[23159] <= 16'hFFFF;
rommem[23160] <= 16'hFFFF;
rommem[23161] <= 16'hFFFF;
rommem[23162] <= 16'hFFFF;
rommem[23163] <= 16'hFFFF;
rommem[23164] <= 16'hFFFF;
rommem[23165] <= 16'hFFFF;
rommem[23166] <= 16'hFFFF;
rommem[23167] <= 16'hFFFF;
rommem[23168] <= 16'hFFFF;
rommem[23169] <= 16'hFFFF;
rommem[23170] <= 16'hFFFF;
rommem[23171] <= 16'hFFFF;
rommem[23172] <= 16'hFFFF;
rommem[23173] <= 16'hFFFF;
rommem[23174] <= 16'hFFFF;
rommem[23175] <= 16'hFFFF;
rommem[23176] <= 16'hFFFF;
rommem[23177] <= 16'hFFFF;
rommem[23178] <= 16'hFFFF;
rommem[23179] <= 16'hFFFF;
rommem[23180] <= 16'hFFFF;
rommem[23181] <= 16'hFFFF;
rommem[23182] <= 16'hFFFF;
rommem[23183] <= 16'hFFFF;
rommem[23184] <= 16'hFFFF;
rommem[23185] <= 16'hFFFF;
rommem[23186] <= 16'hFFFF;
rommem[23187] <= 16'hFFFF;
rommem[23188] <= 16'hFFFF;
rommem[23189] <= 16'hFFFF;
rommem[23190] <= 16'hFFFF;
rommem[23191] <= 16'hFFFF;
rommem[23192] <= 16'hFFFF;
rommem[23193] <= 16'hFFFF;
rommem[23194] <= 16'hFFFF;
rommem[23195] <= 16'hFFFF;
rommem[23196] <= 16'hFFFF;
rommem[23197] <= 16'hFFFF;
rommem[23198] <= 16'hFFFF;
rommem[23199] <= 16'hFFFF;
rommem[23200] <= 16'hFFFF;
rommem[23201] <= 16'hFFFF;
rommem[23202] <= 16'hFFFF;
rommem[23203] <= 16'hFFFF;
rommem[23204] <= 16'hFFFF;
rommem[23205] <= 16'hFFFF;
rommem[23206] <= 16'hFFFF;
rommem[23207] <= 16'hFFFF;
rommem[23208] <= 16'hFFFF;
rommem[23209] <= 16'hFFFF;
rommem[23210] <= 16'hFFFF;
rommem[23211] <= 16'hFFFF;
rommem[23212] <= 16'hFFFF;
rommem[23213] <= 16'hFFFF;
rommem[23214] <= 16'hFFFF;
rommem[23215] <= 16'hFFFF;
rommem[23216] <= 16'hFFFF;
rommem[23217] <= 16'hFFFF;
rommem[23218] <= 16'hFFFF;
rommem[23219] <= 16'hFFFF;
rommem[23220] <= 16'hFFFF;
rommem[23221] <= 16'hFFFF;
rommem[23222] <= 16'hFFFF;
rommem[23223] <= 16'hFFFF;
rommem[23224] <= 16'hFFFF;
rommem[23225] <= 16'hFFFF;
rommem[23226] <= 16'hFFFF;
rommem[23227] <= 16'hFFFF;
rommem[23228] <= 16'hFFFF;
rommem[23229] <= 16'hFFFF;
rommem[23230] <= 16'hFFFF;
rommem[23231] <= 16'hFFFF;
rommem[23232] <= 16'hFFFF;
rommem[23233] <= 16'hFFFF;
rommem[23234] <= 16'hFFFF;
rommem[23235] <= 16'hFFFF;
rommem[23236] <= 16'hFFFF;
rommem[23237] <= 16'hFFFF;
rommem[23238] <= 16'hFFFF;
rommem[23239] <= 16'hFFFF;
rommem[23240] <= 16'hFFFF;
rommem[23241] <= 16'hFFFF;
rommem[23242] <= 16'hFFFF;
rommem[23243] <= 16'hFFFF;
rommem[23244] <= 16'hFFFF;
rommem[23245] <= 16'hFFFF;
rommem[23246] <= 16'hFFFF;
rommem[23247] <= 16'hFFFF;
rommem[23248] <= 16'hFFFF;
rommem[23249] <= 16'hFFFF;
rommem[23250] <= 16'hFFFF;
rommem[23251] <= 16'hFFFF;
rommem[23252] <= 16'hFFFF;
rommem[23253] <= 16'hFFFF;
rommem[23254] <= 16'hFFFF;
rommem[23255] <= 16'hFFFF;
rommem[23256] <= 16'hFFFF;
rommem[23257] <= 16'hFFFF;
rommem[23258] <= 16'hFFFF;
rommem[23259] <= 16'hFFFF;
rommem[23260] <= 16'hFFFF;
rommem[23261] <= 16'hFFFF;
rommem[23262] <= 16'hFFFF;
rommem[23263] <= 16'hFFFF;
rommem[23264] <= 16'hFFFF;
rommem[23265] <= 16'hFFFF;
rommem[23266] <= 16'hFFFF;
rommem[23267] <= 16'hFFFF;
rommem[23268] <= 16'hFFFF;
rommem[23269] <= 16'hFFFF;
rommem[23270] <= 16'hFFFF;
rommem[23271] <= 16'hFFFF;
rommem[23272] <= 16'hFFFF;
rommem[23273] <= 16'hFFFF;
rommem[23274] <= 16'hFFFF;
rommem[23275] <= 16'hFFFF;
rommem[23276] <= 16'hFFFF;
rommem[23277] <= 16'hFFFF;
rommem[23278] <= 16'hFFFF;
rommem[23279] <= 16'hFFFF;
rommem[23280] <= 16'hFFFF;
rommem[23281] <= 16'hFFFF;
rommem[23282] <= 16'hFFFF;
rommem[23283] <= 16'hFFFF;
rommem[23284] <= 16'hFFFF;
rommem[23285] <= 16'hFFFF;
rommem[23286] <= 16'hFFFF;
rommem[23287] <= 16'hFFFF;
rommem[23288] <= 16'hFFFF;
rommem[23289] <= 16'hFFFF;
rommem[23290] <= 16'hFFFF;
rommem[23291] <= 16'hFFFF;
rommem[23292] <= 16'hFFFF;
rommem[23293] <= 16'hFFFF;
rommem[23294] <= 16'hFFFF;
rommem[23295] <= 16'hFFFF;
rommem[23296] <= 16'hFFFF;
rommem[23297] <= 16'hFFFF;
rommem[23298] <= 16'hFFFF;
rommem[23299] <= 16'hFFFF;
rommem[23300] <= 16'hFFFF;
rommem[23301] <= 16'hFFFF;
rommem[23302] <= 16'hFFFF;
rommem[23303] <= 16'hFFFF;
rommem[23304] <= 16'hFFFF;
rommem[23305] <= 16'hFFFF;
rommem[23306] <= 16'hFFFF;
rommem[23307] <= 16'hFFFF;
rommem[23308] <= 16'hFFFF;
rommem[23309] <= 16'hFFFF;
rommem[23310] <= 16'hFFFF;
rommem[23311] <= 16'hFFFF;
rommem[23312] <= 16'hFFFF;
rommem[23313] <= 16'hFFFF;
rommem[23314] <= 16'hFFFF;
rommem[23315] <= 16'hFFFF;
rommem[23316] <= 16'hFFFF;
rommem[23317] <= 16'hFFFF;
rommem[23318] <= 16'hFFFF;
rommem[23319] <= 16'hFFFF;
rommem[23320] <= 16'hFFFF;
rommem[23321] <= 16'hFFFF;
rommem[23322] <= 16'hFFFF;
rommem[23323] <= 16'hFFFF;
rommem[23324] <= 16'hFFFF;
rommem[23325] <= 16'hFFFF;
rommem[23326] <= 16'hFFFF;
rommem[23327] <= 16'hFFFF;
rommem[23328] <= 16'hFFFF;
rommem[23329] <= 16'hFFFF;
rommem[23330] <= 16'hFFFF;
rommem[23331] <= 16'hFFFF;
rommem[23332] <= 16'hFFFF;
rommem[23333] <= 16'hFFFF;
rommem[23334] <= 16'hFFFF;
rommem[23335] <= 16'hFFFF;
rommem[23336] <= 16'hFFFF;
rommem[23337] <= 16'hFFFF;
rommem[23338] <= 16'hFFFF;
rommem[23339] <= 16'hFFFF;
rommem[23340] <= 16'hFFFF;
rommem[23341] <= 16'hFFFF;
rommem[23342] <= 16'hFFFF;
rommem[23343] <= 16'hFFFF;
rommem[23344] <= 16'hFFFF;
rommem[23345] <= 16'hFFFF;
rommem[23346] <= 16'hFFFF;
rommem[23347] <= 16'hFFFF;
rommem[23348] <= 16'hFFFF;
rommem[23349] <= 16'hFFFF;
rommem[23350] <= 16'hFFFF;
rommem[23351] <= 16'hFFFF;
rommem[23352] <= 16'hFFFF;
rommem[23353] <= 16'hFFFF;
rommem[23354] <= 16'hFFFF;
rommem[23355] <= 16'hFFFF;
rommem[23356] <= 16'hFFFF;
rommem[23357] <= 16'hFFFF;
rommem[23358] <= 16'hFFFF;
rommem[23359] <= 16'hFFFF;
rommem[23360] <= 16'hFFFF;
rommem[23361] <= 16'hFFFF;
rommem[23362] <= 16'hFFFF;
rommem[23363] <= 16'hFFFF;
rommem[23364] <= 16'hFFFF;
rommem[23365] <= 16'hFFFF;
rommem[23366] <= 16'hFFFF;
rommem[23367] <= 16'hFFFF;
rommem[23368] <= 16'hFFFF;
rommem[23369] <= 16'hFFFF;
rommem[23370] <= 16'hFFFF;
rommem[23371] <= 16'hFFFF;
rommem[23372] <= 16'hFFFF;
rommem[23373] <= 16'hFFFF;
rommem[23374] <= 16'hFFFF;
rommem[23375] <= 16'hFFFF;
rommem[23376] <= 16'hFFFF;
rommem[23377] <= 16'hFFFF;
rommem[23378] <= 16'hFFFF;
rommem[23379] <= 16'hFFFF;
rommem[23380] <= 16'hFFFF;
rommem[23381] <= 16'hFFFF;
rommem[23382] <= 16'hFFFF;
rommem[23383] <= 16'hFFFF;
rommem[23384] <= 16'hFFFF;
rommem[23385] <= 16'hFFFF;
rommem[23386] <= 16'hFFFF;
rommem[23387] <= 16'hFFFF;
rommem[23388] <= 16'hFFFF;
rommem[23389] <= 16'hFFFF;
rommem[23390] <= 16'hFFFF;
rommem[23391] <= 16'hFFFF;
rommem[23392] <= 16'hFFFF;
rommem[23393] <= 16'hFFFF;
rommem[23394] <= 16'hFFFF;
rommem[23395] <= 16'hFFFF;
rommem[23396] <= 16'hFFFF;
rommem[23397] <= 16'hFFFF;
rommem[23398] <= 16'hFFFF;
rommem[23399] <= 16'hFFFF;
rommem[23400] <= 16'hFFFF;
rommem[23401] <= 16'hFFFF;
rommem[23402] <= 16'hFFFF;
rommem[23403] <= 16'hFFFF;
rommem[23404] <= 16'hFFFF;
rommem[23405] <= 16'hFFFF;
rommem[23406] <= 16'hFFFF;
rommem[23407] <= 16'hFFFF;
rommem[23408] <= 16'hFFFF;
rommem[23409] <= 16'hFFFF;
rommem[23410] <= 16'hFFFF;
rommem[23411] <= 16'hFFFF;
rommem[23412] <= 16'hFFFF;
rommem[23413] <= 16'hFFFF;
rommem[23414] <= 16'hFFFF;
rommem[23415] <= 16'hFFFF;
rommem[23416] <= 16'hFFFF;
rommem[23417] <= 16'hFFFF;
rommem[23418] <= 16'hFFFF;
rommem[23419] <= 16'hFFFF;
rommem[23420] <= 16'hFFFF;
rommem[23421] <= 16'hFFFF;
rommem[23422] <= 16'hFFFF;
rommem[23423] <= 16'hFFFF;
rommem[23424] <= 16'hFFFF;
rommem[23425] <= 16'hFFFF;
rommem[23426] <= 16'hFFFF;
rommem[23427] <= 16'hFFFF;
rommem[23428] <= 16'hFFFF;
rommem[23429] <= 16'hFFFF;
rommem[23430] <= 16'hFFFF;
rommem[23431] <= 16'hFFFF;
rommem[23432] <= 16'hFFFF;
rommem[23433] <= 16'hFFFF;
rommem[23434] <= 16'hFFFF;
rommem[23435] <= 16'hFFFF;
rommem[23436] <= 16'hFFFF;
rommem[23437] <= 16'hFFFF;
rommem[23438] <= 16'hFFFF;
rommem[23439] <= 16'hFFFF;
rommem[23440] <= 16'hFFFF;
rommem[23441] <= 16'hFFFF;
rommem[23442] <= 16'hFFFF;
rommem[23443] <= 16'hFFFF;
rommem[23444] <= 16'hFFFF;
rommem[23445] <= 16'hFFFF;
rommem[23446] <= 16'hFFFF;
rommem[23447] <= 16'hFFFF;
rommem[23448] <= 16'hFFFF;
rommem[23449] <= 16'hFFFF;
rommem[23450] <= 16'hFFFF;
rommem[23451] <= 16'hFFFF;
rommem[23452] <= 16'hFFFF;
rommem[23453] <= 16'hFFFF;
rommem[23454] <= 16'hFFFF;
rommem[23455] <= 16'hFFFF;
rommem[23456] <= 16'hFFFF;
rommem[23457] <= 16'hFFFF;
rommem[23458] <= 16'hFFFF;
rommem[23459] <= 16'hFFFF;
rommem[23460] <= 16'hFFFF;
rommem[23461] <= 16'hFFFF;
rommem[23462] <= 16'hFFFF;
rommem[23463] <= 16'hFFFF;
rommem[23464] <= 16'hFFFF;
rommem[23465] <= 16'hFFFF;
rommem[23466] <= 16'hFFFF;
rommem[23467] <= 16'hFFFF;
rommem[23468] <= 16'hFFFF;
rommem[23469] <= 16'hFFFF;
rommem[23470] <= 16'hFFFF;
rommem[23471] <= 16'hFFFF;
rommem[23472] <= 16'hFFFF;
rommem[23473] <= 16'hFFFF;
rommem[23474] <= 16'hFFFF;
rommem[23475] <= 16'hFFFF;
rommem[23476] <= 16'hFFFF;
rommem[23477] <= 16'hFFFF;
rommem[23478] <= 16'hFFFF;
rommem[23479] <= 16'hFFFF;
rommem[23480] <= 16'hFFFF;
rommem[23481] <= 16'hFFFF;
rommem[23482] <= 16'hFFFF;
rommem[23483] <= 16'hFFFF;
rommem[23484] <= 16'hFFFF;
rommem[23485] <= 16'hFFFF;
rommem[23486] <= 16'hFFFF;
rommem[23487] <= 16'hFFFF;
rommem[23488] <= 16'hFFFF;
rommem[23489] <= 16'hFFFF;
rommem[23490] <= 16'hFFFF;
rommem[23491] <= 16'hFFFF;
rommem[23492] <= 16'hFFFF;
rommem[23493] <= 16'hFFFF;
rommem[23494] <= 16'hFFFF;
rommem[23495] <= 16'hFFFF;
rommem[23496] <= 16'hFFFF;
rommem[23497] <= 16'hFFFF;
rommem[23498] <= 16'hFFFF;
rommem[23499] <= 16'hFFFF;
rommem[23500] <= 16'hFFFF;
rommem[23501] <= 16'hFFFF;
rommem[23502] <= 16'hFFFF;
rommem[23503] <= 16'hFFFF;
rommem[23504] <= 16'hFFFF;
rommem[23505] <= 16'hFFFF;
rommem[23506] <= 16'hFFFF;
rommem[23507] <= 16'hFFFF;
rommem[23508] <= 16'hFFFF;
rommem[23509] <= 16'hFFFF;
rommem[23510] <= 16'hFFFF;
rommem[23511] <= 16'hFFFF;
rommem[23512] <= 16'hFFFF;
rommem[23513] <= 16'hFFFF;
rommem[23514] <= 16'hFFFF;
rommem[23515] <= 16'hFFFF;
rommem[23516] <= 16'hFFFF;
rommem[23517] <= 16'hFFFF;
rommem[23518] <= 16'hFFFF;
rommem[23519] <= 16'hFFFF;
rommem[23520] <= 16'hFFFF;
rommem[23521] <= 16'hFFFF;
rommem[23522] <= 16'hFFFF;
rommem[23523] <= 16'hFFFF;
rommem[23524] <= 16'hFFFF;
rommem[23525] <= 16'hFFFF;
rommem[23526] <= 16'hFFFF;
rommem[23527] <= 16'hFFFF;
rommem[23528] <= 16'hFFFF;
rommem[23529] <= 16'hFFFF;
rommem[23530] <= 16'hFFFF;
rommem[23531] <= 16'hFFFF;
rommem[23532] <= 16'hFFFF;
rommem[23533] <= 16'hFFFF;
rommem[23534] <= 16'hFFFF;
rommem[23535] <= 16'hFFFF;
rommem[23536] <= 16'hFFFF;
rommem[23537] <= 16'hFFFF;
rommem[23538] <= 16'hFFFF;
rommem[23539] <= 16'hFFFF;
rommem[23540] <= 16'hFFFF;
rommem[23541] <= 16'hFFFF;
rommem[23542] <= 16'hFFFF;
rommem[23543] <= 16'hFFFF;
rommem[23544] <= 16'hFFFF;
rommem[23545] <= 16'hFFFF;
rommem[23546] <= 16'hFFFF;
rommem[23547] <= 16'hFFFF;
rommem[23548] <= 16'hFFFF;
rommem[23549] <= 16'hFFFF;
rommem[23550] <= 16'hFFFF;
rommem[23551] <= 16'hFFFF;
rommem[23552] <= 16'hFFFF;
rommem[23553] <= 16'hFFFF;
rommem[23554] <= 16'hFFFF;
rommem[23555] <= 16'hFFFF;
rommem[23556] <= 16'hFFFF;
rommem[23557] <= 16'hFFFF;
rommem[23558] <= 16'hFFFF;
rommem[23559] <= 16'hFFFF;
rommem[23560] <= 16'hFFFF;
rommem[23561] <= 16'hFFFF;
rommem[23562] <= 16'hFFFF;
rommem[23563] <= 16'hFFFF;
rommem[23564] <= 16'hFFFF;
rommem[23565] <= 16'hFFFF;
rommem[23566] <= 16'hFFFF;
rommem[23567] <= 16'hFFFF;
rommem[23568] <= 16'hFFFF;
rommem[23569] <= 16'hFFFF;
rommem[23570] <= 16'hFFFF;
rommem[23571] <= 16'hFFFF;
rommem[23572] <= 16'hFFFF;
rommem[23573] <= 16'hFFFF;
rommem[23574] <= 16'hFFFF;
rommem[23575] <= 16'hFFFF;
rommem[23576] <= 16'hFFFF;
rommem[23577] <= 16'hFFFF;
rommem[23578] <= 16'hFFFF;
rommem[23579] <= 16'hFFFF;
rommem[23580] <= 16'hFFFF;
rommem[23581] <= 16'hFFFF;
rommem[23582] <= 16'hFFFF;
rommem[23583] <= 16'hFFFF;
rommem[23584] <= 16'hFFFF;
rommem[23585] <= 16'hFFFF;
rommem[23586] <= 16'hFFFF;
rommem[23587] <= 16'hFFFF;
rommem[23588] <= 16'hFFFF;
rommem[23589] <= 16'hFFFF;
rommem[23590] <= 16'hFFFF;
rommem[23591] <= 16'hFFFF;
rommem[23592] <= 16'hFFFF;
rommem[23593] <= 16'hFFFF;
rommem[23594] <= 16'hFFFF;
rommem[23595] <= 16'hFFFF;
rommem[23596] <= 16'hFFFF;
rommem[23597] <= 16'hFFFF;
rommem[23598] <= 16'hFFFF;
rommem[23599] <= 16'hFFFF;
rommem[23600] <= 16'hFFFF;
rommem[23601] <= 16'hFFFF;
rommem[23602] <= 16'hFFFF;
rommem[23603] <= 16'hFFFF;
rommem[23604] <= 16'hFFFF;
rommem[23605] <= 16'hFFFF;
rommem[23606] <= 16'hFFFF;
rommem[23607] <= 16'hFFFF;
rommem[23608] <= 16'hFFFF;
rommem[23609] <= 16'hFFFF;
rommem[23610] <= 16'hFFFF;
rommem[23611] <= 16'hFFFF;
rommem[23612] <= 16'hFFFF;
rommem[23613] <= 16'hFFFF;
rommem[23614] <= 16'hFFFF;
rommem[23615] <= 16'hFFFF;
rommem[23616] <= 16'hFFFF;
rommem[23617] <= 16'hFFFF;
rommem[23618] <= 16'hFFFF;
rommem[23619] <= 16'hFFFF;
rommem[23620] <= 16'hFFFF;
rommem[23621] <= 16'hFFFF;
rommem[23622] <= 16'hFFFF;
rommem[23623] <= 16'hFFFF;
rommem[23624] <= 16'hFFFF;
rommem[23625] <= 16'hFFFF;
rommem[23626] <= 16'hFFFF;
rommem[23627] <= 16'hFFFF;
rommem[23628] <= 16'hFFFF;
rommem[23629] <= 16'hFFFF;
rommem[23630] <= 16'hFFFF;
rommem[23631] <= 16'hFFFF;
rommem[23632] <= 16'hFFFF;
rommem[23633] <= 16'hFFFF;
rommem[23634] <= 16'hFFFF;
rommem[23635] <= 16'hFFFF;
rommem[23636] <= 16'hFFFF;
rommem[23637] <= 16'hFFFF;
rommem[23638] <= 16'hFFFF;
rommem[23639] <= 16'hFFFF;
rommem[23640] <= 16'hFFFF;
rommem[23641] <= 16'hFFFF;
rommem[23642] <= 16'hFFFF;
rommem[23643] <= 16'hFFFF;
rommem[23644] <= 16'hFFFF;
rommem[23645] <= 16'hFFFF;
rommem[23646] <= 16'hFFFF;
rommem[23647] <= 16'hFFFF;
rommem[23648] <= 16'hFFFF;
rommem[23649] <= 16'hFFFF;
rommem[23650] <= 16'hFFFF;
rommem[23651] <= 16'hFFFF;
rommem[23652] <= 16'hFFFF;
rommem[23653] <= 16'hFFFF;
rommem[23654] <= 16'hFFFF;
rommem[23655] <= 16'hFFFF;
rommem[23656] <= 16'hFFFF;
rommem[23657] <= 16'hFFFF;
rommem[23658] <= 16'hFFFF;
rommem[23659] <= 16'hFFFF;
rommem[23660] <= 16'hFFFF;
rommem[23661] <= 16'hFFFF;
rommem[23662] <= 16'hFFFF;
rommem[23663] <= 16'hFFFF;
rommem[23664] <= 16'hFFFF;
rommem[23665] <= 16'hFFFF;
rommem[23666] <= 16'hFFFF;
rommem[23667] <= 16'hFFFF;
rommem[23668] <= 16'hFFFF;
rommem[23669] <= 16'hFFFF;
rommem[23670] <= 16'hFFFF;
rommem[23671] <= 16'hFFFF;
rommem[23672] <= 16'hFFFF;
rommem[23673] <= 16'hFFFF;
rommem[23674] <= 16'hFFFF;
rommem[23675] <= 16'hFFFF;
rommem[23676] <= 16'hFFFF;
rommem[23677] <= 16'hFFFF;
rommem[23678] <= 16'hFFFF;
rommem[23679] <= 16'hFFFF;
rommem[23680] <= 16'hFFFF;
rommem[23681] <= 16'hFFFF;
rommem[23682] <= 16'hFFFF;
rommem[23683] <= 16'hFFFF;
rommem[23684] <= 16'hFFFF;
rommem[23685] <= 16'hFFFF;
rommem[23686] <= 16'hFFFF;
rommem[23687] <= 16'hFFFF;
rommem[23688] <= 16'hFFFF;
rommem[23689] <= 16'hFFFF;
rommem[23690] <= 16'hFFFF;
rommem[23691] <= 16'hFFFF;
rommem[23692] <= 16'hFFFF;
rommem[23693] <= 16'hFFFF;
rommem[23694] <= 16'hFFFF;
rommem[23695] <= 16'hFFFF;
rommem[23696] <= 16'hFFFF;
rommem[23697] <= 16'hFFFF;
rommem[23698] <= 16'hFFFF;
rommem[23699] <= 16'hFFFF;
rommem[23700] <= 16'hFFFF;
rommem[23701] <= 16'hFFFF;
rommem[23702] <= 16'hFFFF;
rommem[23703] <= 16'hFFFF;
rommem[23704] <= 16'hFFFF;
rommem[23705] <= 16'hFFFF;
rommem[23706] <= 16'hFFFF;
rommem[23707] <= 16'hFFFF;
rommem[23708] <= 16'hFFFF;
rommem[23709] <= 16'hFFFF;
rommem[23710] <= 16'hFFFF;
rommem[23711] <= 16'hFFFF;
rommem[23712] <= 16'hFFFF;
rommem[23713] <= 16'hFFFF;
rommem[23714] <= 16'hFFFF;
rommem[23715] <= 16'hFFFF;
rommem[23716] <= 16'hFFFF;
rommem[23717] <= 16'hFFFF;
rommem[23718] <= 16'hFFFF;
rommem[23719] <= 16'hFFFF;
rommem[23720] <= 16'hFFFF;
rommem[23721] <= 16'hFFFF;
rommem[23722] <= 16'hFFFF;
rommem[23723] <= 16'hFFFF;
rommem[23724] <= 16'hFFFF;
rommem[23725] <= 16'hFFFF;
rommem[23726] <= 16'hFFFF;
rommem[23727] <= 16'hFFFF;
rommem[23728] <= 16'hFFFF;
rommem[23729] <= 16'hFFFF;
rommem[23730] <= 16'hFFFF;
rommem[23731] <= 16'hFFFF;
rommem[23732] <= 16'hFFFF;
rommem[23733] <= 16'hFFFF;
rommem[23734] <= 16'hFFFF;
rommem[23735] <= 16'hFFFF;
rommem[23736] <= 16'hFFFF;
rommem[23737] <= 16'hFFFF;
rommem[23738] <= 16'hFFFF;
rommem[23739] <= 16'hFFFF;
rommem[23740] <= 16'hFFFF;
rommem[23741] <= 16'hFFFF;
rommem[23742] <= 16'hFFFF;
rommem[23743] <= 16'hFFFF;
rommem[23744] <= 16'hFFFF;
rommem[23745] <= 16'hFFFF;
rommem[23746] <= 16'hFFFF;
rommem[23747] <= 16'hFFFF;
rommem[23748] <= 16'hFFFF;
rommem[23749] <= 16'hFFFF;
rommem[23750] <= 16'hFFFF;
rommem[23751] <= 16'hFFFF;
rommem[23752] <= 16'hFFFF;
rommem[23753] <= 16'hFFFF;
rommem[23754] <= 16'hFFFF;
rommem[23755] <= 16'hFFFF;
rommem[23756] <= 16'hFFFF;
rommem[23757] <= 16'hFFFF;
rommem[23758] <= 16'hFFFF;
rommem[23759] <= 16'hFFFF;
rommem[23760] <= 16'hFFFF;
rommem[23761] <= 16'hFFFF;
rommem[23762] <= 16'hFFFF;
rommem[23763] <= 16'hFFFF;
rommem[23764] <= 16'hFFFF;
rommem[23765] <= 16'hFFFF;
rommem[23766] <= 16'hFFFF;
rommem[23767] <= 16'hFFFF;
rommem[23768] <= 16'hFFFF;
rommem[23769] <= 16'hFFFF;
rommem[23770] <= 16'hFFFF;
rommem[23771] <= 16'hFFFF;
rommem[23772] <= 16'hFFFF;
rommem[23773] <= 16'hFFFF;
rommem[23774] <= 16'hFFFF;
rommem[23775] <= 16'hFFFF;
rommem[23776] <= 16'hFFFF;
rommem[23777] <= 16'hFFFF;
rommem[23778] <= 16'hFFFF;
rommem[23779] <= 16'hFFFF;
rommem[23780] <= 16'hFFFF;
rommem[23781] <= 16'hFFFF;
rommem[23782] <= 16'hFFFF;
rommem[23783] <= 16'hFFFF;
rommem[23784] <= 16'hFFFF;
rommem[23785] <= 16'hFFFF;
rommem[23786] <= 16'hFFFF;
rommem[23787] <= 16'hFFFF;
rommem[23788] <= 16'hFFFF;
rommem[23789] <= 16'hFFFF;
rommem[23790] <= 16'hFFFF;
rommem[23791] <= 16'hFFFF;
rommem[23792] <= 16'hFFFF;
rommem[23793] <= 16'hFFFF;
rommem[23794] <= 16'hFFFF;
rommem[23795] <= 16'hFFFF;
rommem[23796] <= 16'hFFFF;
rommem[23797] <= 16'hFFFF;
rommem[23798] <= 16'hFFFF;
rommem[23799] <= 16'hFFFF;
rommem[23800] <= 16'hFFFF;
rommem[23801] <= 16'hFFFF;
rommem[23802] <= 16'hFFFF;
rommem[23803] <= 16'hFFFF;
rommem[23804] <= 16'hFFFF;
rommem[23805] <= 16'hFFFF;
rommem[23806] <= 16'hFFFF;
rommem[23807] <= 16'hFFFF;
rommem[23808] <= 16'hFFFF;
rommem[23809] <= 16'hFFFF;
rommem[23810] <= 16'hFFFF;
rommem[23811] <= 16'hFFFF;
rommem[23812] <= 16'hFFFF;
rommem[23813] <= 16'hFFFF;
rommem[23814] <= 16'hFFFF;
rommem[23815] <= 16'hFFFF;
rommem[23816] <= 16'hFFFF;
rommem[23817] <= 16'hFFFF;
rommem[23818] <= 16'hFFFF;
rommem[23819] <= 16'hFFFF;
rommem[23820] <= 16'hFFFF;
rommem[23821] <= 16'hFFFF;
rommem[23822] <= 16'hFFFF;
rommem[23823] <= 16'hFFFF;
rommem[23824] <= 16'hFFFF;
rommem[23825] <= 16'hFFFF;
rommem[23826] <= 16'hFFFF;
rommem[23827] <= 16'hFFFF;
rommem[23828] <= 16'hFFFF;
rommem[23829] <= 16'hFFFF;
rommem[23830] <= 16'hFFFF;
rommem[23831] <= 16'hFFFF;
rommem[23832] <= 16'hFFFF;
rommem[23833] <= 16'hFFFF;
rommem[23834] <= 16'hFFFF;
rommem[23835] <= 16'hFFFF;
rommem[23836] <= 16'hFFFF;
rommem[23837] <= 16'hFFFF;
rommem[23838] <= 16'hFFFF;
rommem[23839] <= 16'hFFFF;
rommem[23840] <= 16'hFFFF;
rommem[23841] <= 16'hFFFF;
rommem[23842] <= 16'hFFFF;
rommem[23843] <= 16'hFFFF;
rommem[23844] <= 16'hFFFF;
rommem[23845] <= 16'hFFFF;
rommem[23846] <= 16'hFFFF;
rommem[23847] <= 16'hFFFF;
rommem[23848] <= 16'hFFFF;
rommem[23849] <= 16'hFFFF;
rommem[23850] <= 16'hFFFF;
rommem[23851] <= 16'hFFFF;
rommem[23852] <= 16'hFFFF;
rommem[23853] <= 16'hFFFF;
rommem[23854] <= 16'hFFFF;
rommem[23855] <= 16'hFFFF;
rommem[23856] <= 16'hFFFF;
rommem[23857] <= 16'hFFFF;
rommem[23858] <= 16'hFFFF;
rommem[23859] <= 16'hFFFF;
rommem[23860] <= 16'hFFFF;
rommem[23861] <= 16'hFFFF;
rommem[23862] <= 16'hFFFF;
rommem[23863] <= 16'hFFFF;
rommem[23864] <= 16'hFFFF;
rommem[23865] <= 16'hFFFF;
rommem[23866] <= 16'hFFFF;
rommem[23867] <= 16'hFFFF;
rommem[23868] <= 16'hFFFF;
rommem[23869] <= 16'hFFFF;
rommem[23870] <= 16'hFFFF;
rommem[23871] <= 16'hFFFF;
rommem[23872] <= 16'hFFFF;
rommem[23873] <= 16'hFFFF;
rommem[23874] <= 16'hFFFF;
rommem[23875] <= 16'hFFFF;
rommem[23876] <= 16'hFFFF;
rommem[23877] <= 16'hFFFF;
rommem[23878] <= 16'hFFFF;
rommem[23879] <= 16'hFFFF;
rommem[23880] <= 16'hFFFF;
rommem[23881] <= 16'hFFFF;
rommem[23882] <= 16'hFFFF;
rommem[23883] <= 16'hFFFF;
rommem[23884] <= 16'hFFFF;
rommem[23885] <= 16'hFFFF;
rommem[23886] <= 16'hFFFF;
rommem[23887] <= 16'hFFFF;
rommem[23888] <= 16'hFFFF;
rommem[23889] <= 16'hFFFF;
rommem[23890] <= 16'hFFFF;
rommem[23891] <= 16'hFFFF;
rommem[23892] <= 16'hFFFF;
rommem[23893] <= 16'hFFFF;
rommem[23894] <= 16'hFFFF;
rommem[23895] <= 16'hFFFF;
rommem[23896] <= 16'hFFFF;
rommem[23897] <= 16'hFFFF;
rommem[23898] <= 16'hFFFF;
rommem[23899] <= 16'hFFFF;
rommem[23900] <= 16'hFFFF;
rommem[23901] <= 16'hFFFF;
rommem[23902] <= 16'hFFFF;
rommem[23903] <= 16'hFFFF;
rommem[23904] <= 16'hFFFF;
rommem[23905] <= 16'hFFFF;
rommem[23906] <= 16'hFFFF;
rommem[23907] <= 16'hFFFF;
rommem[23908] <= 16'hFFFF;
rommem[23909] <= 16'hFFFF;
rommem[23910] <= 16'hFFFF;
rommem[23911] <= 16'hFFFF;
rommem[23912] <= 16'hFFFF;
rommem[23913] <= 16'hFFFF;
rommem[23914] <= 16'hFFFF;
rommem[23915] <= 16'hFFFF;
rommem[23916] <= 16'hFFFF;
rommem[23917] <= 16'hFFFF;
rommem[23918] <= 16'hFFFF;
rommem[23919] <= 16'hFFFF;
rommem[23920] <= 16'hFFFF;
rommem[23921] <= 16'hFFFF;
rommem[23922] <= 16'hFFFF;
rommem[23923] <= 16'hFFFF;
rommem[23924] <= 16'hFFFF;
rommem[23925] <= 16'hFFFF;
rommem[23926] <= 16'hFFFF;
rommem[23927] <= 16'hFFFF;
rommem[23928] <= 16'hFFFF;
rommem[23929] <= 16'hFFFF;
rommem[23930] <= 16'hFFFF;
rommem[23931] <= 16'hFFFF;
rommem[23932] <= 16'hFFFF;
rommem[23933] <= 16'hFFFF;
rommem[23934] <= 16'hFFFF;
rommem[23935] <= 16'hFFFF;
rommem[23936] <= 16'hFFFF;
rommem[23937] <= 16'hFFFF;
rommem[23938] <= 16'hFFFF;
rommem[23939] <= 16'hFFFF;
rommem[23940] <= 16'hFFFF;
rommem[23941] <= 16'hFFFF;
rommem[23942] <= 16'hFFFF;
rommem[23943] <= 16'hFFFF;
rommem[23944] <= 16'hFFFF;
rommem[23945] <= 16'hFFFF;
rommem[23946] <= 16'hFFFF;
rommem[23947] <= 16'hFFFF;
rommem[23948] <= 16'hFFFF;
rommem[23949] <= 16'hFFFF;
rommem[23950] <= 16'hFFFF;
rommem[23951] <= 16'hFFFF;
rommem[23952] <= 16'hFFFF;
rommem[23953] <= 16'hFFFF;
rommem[23954] <= 16'hFFFF;
rommem[23955] <= 16'hFFFF;
rommem[23956] <= 16'hFFFF;
rommem[23957] <= 16'hFFFF;
rommem[23958] <= 16'hFFFF;
rommem[23959] <= 16'hFFFF;
rommem[23960] <= 16'hFFFF;
rommem[23961] <= 16'hFFFF;
rommem[23962] <= 16'hFFFF;
rommem[23963] <= 16'hFFFF;
rommem[23964] <= 16'hFFFF;
rommem[23965] <= 16'hFFFF;
rommem[23966] <= 16'hFFFF;
rommem[23967] <= 16'hFFFF;
rommem[23968] <= 16'hFFFF;
rommem[23969] <= 16'hFFFF;
rommem[23970] <= 16'hFFFF;
rommem[23971] <= 16'hFFFF;
rommem[23972] <= 16'hFFFF;
rommem[23973] <= 16'hFFFF;
rommem[23974] <= 16'hFFFF;
rommem[23975] <= 16'hFFFF;
rommem[23976] <= 16'hFFFF;
rommem[23977] <= 16'hFFFF;
rommem[23978] <= 16'hFFFF;
rommem[23979] <= 16'hFFFF;
rommem[23980] <= 16'hFFFF;
rommem[23981] <= 16'hFFFF;
rommem[23982] <= 16'hFFFF;
rommem[23983] <= 16'hFFFF;
rommem[23984] <= 16'hFFFF;
rommem[23985] <= 16'hFFFF;
rommem[23986] <= 16'hFFFF;
rommem[23987] <= 16'hFFFF;
rommem[23988] <= 16'hFFFF;
rommem[23989] <= 16'hFFFF;
rommem[23990] <= 16'hFFFF;
rommem[23991] <= 16'hFFFF;
rommem[23992] <= 16'hFFFF;
rommem[23993] <= 16'hFFFF;
rommem[23994] <= 16'hFFFF;
rommem[23995] <= 16'hFFFF;
rommem[23996] <= 16'hFFFF;
rommem[23997] <= 16'hFFFF;
rommem[23998] <= 16'hFFFF;
rommem[23999] <= 16'hFFFF;
rommem[24000] <= 16'hFFFF;
rommem[24001] <= 16'hFFFF;
rommem[24002] <= 16'hFFFF;
rommem[24003] <= 16'hFFFF;
rommem[24004] <= 16'hFFFF;
rommem[24005] <= 16'hFFFF;
rommem[24006] <= 16'hFFFF;
rommem[24007] <= 16'hFFFF;
rommem[24008] <= 16'hFFFF;
rommem[24009] <= 16'hFFFF;
rommem[24010] <= 16'hFFFF;
rommem[24011] <= 16'hFFFF;
rommem[24012] <= 16'hFFFF;
rommem[24013] <= 16'hFFFF;
rommem[24014] <= 16'hFFFF;
rommem[24015] <= 16'hFFFF;
rommem[24016] <= 16'hFFFF;
rommem[24017] <= 16'hFFFF;
rommem[24018] <= 16'hFFFF;
rommem[24019] <= 16'hFFFF;
rommem[24020] <= 16'hFFFF;
rommem[24021] <= 16'hFFFF;
rommem[24022] <= 16'hFFFF;
rommem[24023] <= 16'hFFFF;
rommem[24024] <= 16'hFFFF;
rommem[24025] <= 16'hFFFF;
rommem[24026] <= 16'hFFFF;
rommem[24027] <= 16'hFFFF;
rommem[24028] <= 16'hFFFF;
rommem[24029] <= 16'hFFFF;
rommem[24030] <= 16'hFFFF;
rommem[24031] <= 16'hFFFF;
rommem[24032] <= 16'hFFFF;
rommem[24033] <= 16'hFFFF;
rommem[24034] <= 16'hFFFF;
rommem[24035] <= 16'hFFFF;
rommem[24036] <= 16'hFFFF;
rommem[24037] <= 16'hFFFF;
rommem[24038] <= 16'hFFFF;
rommem[24039] <= 16'hFFFF;
rommem[24040] <= 16'hFFFF;
rommem[24041] <= 16'hFFFF;
rommem[24042] <= 16'hFFFF;
rommem[24043] <= 16'hFFFF;
rommem[24044] <= 16'hFFFF;
rommem[24045] <= 16'hFFFF;
rommem[24046] <= 16'hFFFF;
rommem[24047] <= 16'hFFFF;
rommem[24048] <= 16'hFFFF;
rommem[24049] <= 16'hFFFF;
rommem[24050] <= 16'hFFFF;
rommem[24051] <= 16'hFFFF;
rommem[24052] <= 16'hFFFF;
rommem[24053] <= 16'hFFFF;
rommem[24054] <= 16'hFFFF;
rommem[24055] <= 16'hFFFF;
rommem[24056] <= 16'hFFFF;
rommem[24057] <= 16'hFFFF;
rommem[24058] <= 16'hFFFF;
rommem[24059] <= 16'hFFFF;
rommem[24060] <= 16'hFFFF;
rommem[24061] <= 16'hFFFF;
rommem[24062] <= 16'hFFFF;
rommem[24063] <= 16'hFFFF;
rommem[24064] <= 16'hFFFF;
rommem[24065] <= 16'hFFFF;
rommem[24066] <= 16'hFFFF;
rommem[24067] <= 16'hFFFF;
rommem[24068] <= 16'hFFFF;
rommem[24069] <= 16'hFFFF;
rommem[24070] <= 16'hFFFF;
rommem[24071] <= 16'hFFFF;
rommem[24072] <= 16'hFFFF;
rommem[24073] <= 16'hFFFF;
rommem[24074] <= 16'hFFFF;
rommem[24075] <= 16'hFFFF;
rommem[24076] <= 16'hFFFF;
rommem[24077] <= 16'hFFFF;
rommem[24078] <= 16'hFFFF;
rommem[24079] <= 16'hFFFF;
rommem[24080] <= 16'hFFFF;
rommem[24081] <= 16'hFFFF;
rommem[24082] <= 16'hFFFF;
rommem[24083] <= 16'hFFFF;
rommem[24084] <= 16'hFFFF;
rommem[24085] <= 16'hFFFF;
rommem[24086] <= 16'hFFFF;
rommem[24087] <= 16'hFFFF;
rommem[24088] <= 16'hFFFF;
rommem[24089] <= 16'hFFFF;
rommem[24090] <= 16'hFFFF;
rommem[24091] <= 16'hFFFF;
rommem[24092] <= 16'hFFFF;
rommem[24093] <= 16'hFFFF;
rommem[24094] <= 16'hFFFF;
rommem[24095] <= 16'hFFFF;
rommem[24096] <= 16'hFFFF;
rommem[24097] <= 16'hFFFF;
rommem[24098] <= 16'hFFFF;
rommem[24099] <= 16'hFFFF;
rommem[24100] <= 16'hFFFF;
rommem[24101] <= 16'hFFFF;
rommem[24102] <= 16'hFFFF;
rommem[24103] <= 16'hFFFF;
rommem[24104] <= 16'hFFFF;
rommem[24105] <= 16'hFFFF;
rommem[24106] <= 16'hFFFF;
rommem[24107] <= 16'hFFFF;
rommem[24108] <= 16'hFFFF;
rommem[24109] <= 16'hFFFF;
rommem[24110] <= 16'hFFFF;
rommem[24111] <= 16'hFFFF;
rommem[24112] <= 16'hFFFF;
rommem[24113] <= 16'hFFFF;
rommem[24114] <= 16'hFFFF;
rommem[24115] <= 16'hFFFF;
rommem[24116] <= 16'hFFFF;
rommem[24117] <= 16'hFFFF;
rommem[24118] <= 16'hFFFF;
rommem[24119] <= 16'hFFFF;
rommem[24120] <= 16'hFFFF;
rommem[24121] <= 16'hFFFF;
rommem[24122] <= 16'hFFFF;
rommem[24123] <= 16'hFFFF;
rommem[24124] <= 16'hFFFF;
rommem[24125] <= 16'hFFFF;
rommem[24126] <= 16'hFFFF;
rommem[24127] <= 16'hFFFF;
rommem[24128] <= 16'hFFFF;
rommem[24129] <= 16'hFFFF;
rommem[24130] <= 16'hFFFF;
rommem[24131] <= 16'hFFFF;
rommem[24132] <= 16'hFFFF;
rommem[24133] <= 16'hFFFF;
rommem[24134] <= 16'hFFFF;
rommem[24135] <= 16'hFFFF;
rommem[24136] <= 16'hFFFF;
rommem[24137] <= 16'hFFFF;
rommem[24138] <= 16'hFFFF;
rommem[24139] <= 16'hFFFF;
rommem[24140] <= 16'hFFFF;
rommem[24141] <= 16'hFFFF;
rommem[24142] <= 16'hFFFF;
rommem[24143] <= 16'hFFFF;
rommem[24144] <= 16'hFFFF;
rommem[24145] <= 16'hFFFF;
rommem[24146] <= 16'hFFFF;
rommem[24147] <= 16'hFFFF;
rommem[24148] <= 16'hFFFF;
rommem[24149] <= 16'hFFFF;
rommem[24150] <= 16'hFFFF;
rommem[24151] <= 16'hFFFF;
rommem[24152] <= 16'hFFFF;
rommem[24153] <= 16'hFFFF;
rommem[24154] <= 16'hFFFF;
rommem[24155] <= 16'hFFFF;
rommem[24156] <= 16'hFFFF;
rommem[24157] <= 16'hFFFF;
rommem[24158] <= 16'hFFFF;
rommem[24159] <= 16'hFFFF;
rommem[24160] <= 16'hFFFF;
rommem[24161] <= 16'hFFFF;
rommem[24162] <= 16'hFFFF;
rommem[24163] <= 16'hFFFF;
rommem[24164] <= 16'hFFFF;
rommem[24165] <= 16'hFFFF;
rommem[24166] <= 16'hFFFF;
rommem[24167] <= 16'hFFFF;
rommem[24168] <= 16'hFFFF;
rommem[24169] <= 16'hFFFF;
rommem[24170] <= 16'hFFFF;
rommem[24171] <= 16'hFFFF;
rommem[24172] <= 16'hFFFF;
rommem[24173] <= 16'hFFFF;
rommem[24174] <= 16'hFFFF;
rommem[24175] <= 16'hFFFF;
rommem[24176] <= 16'hFFFF;
rommem[24177] <= 16'hFFFF;
rommem[24178] <= 16'hFFFF;
rommem[24179] <= 16'hFFFF;
rommem[24180] <= 16'hFFFF;
rommem[24181] <= 16'hFFFF;
rommem[24182] <= 16'hFFFF;
rommem[24183] <= 16'hFFFF;
rommem[24184] <= 16'hFFFF;
rommem[24185] <= 16'hFFFF;
rommem[24186] <= 16'hFFFF;
rommem[24187] <= 16'hFFFF;
rommem[24188] <= 16'hFFFF;
rommem[24189] <= 16'hFFFF;
rommem[24190] <= 16'hFFFF;
rommem[24191] <= 16'hFFFF;
rommem[24192] <= 16'hFFFF;
rommem[24193] <= 16'hFFFF;
rommem[24194] <= 16'hFFFF;
rommem[24195] <= 16'hFFFF;
rommem[24196] <= 16'hFFFF;
rommem[24197] <= 16'hFFFF;
rommem[24198] <= 16'hFFFF;
rommem[24199] <= 16'hFFFF;
rommem[24200] <= 16'hFFFF;
rommem[24201] <= 16'hFFFF;
rommem[24202] <= 16'hFFFF;
rommem[24203] <= 16'hFFFF;
rommem[24204] <= 16'hFFFF;
rommem[24205] <= 16'hFFFF;
rommem[24206] <= 16'hFFFF;
rommem[24207] <= 16'hFFFF;
rommem[24208] <= 16'hFFFF;
rommem[24209] <= 16'hFFFF;
rommem[24210] <= 16'hFFFF;
rommem[24211] <= 16'hFFFF;
rommem[24212] <= 16'hFFFF;
rommem[24213] <= 16'hFFFF;
rommem[24214] <= 16'hFFFF;
rommem[24215] <= 16'hFFFF;
rommem[24216] <= 16'hFFFF;
rommem[24217] <= 16'hFFFF;
rommem[24218] <= 16'hFFFF;
rommem[24219] <= 16'hFFFF;
rommem[24220] <= 16'hFFFF;
rommem[24221] <= 16'hFFFF;
rommem[24222] <= 16'hFFFF;
rommem[24223] <= 16'hFFFF;
rommem[24224] <= 16'hFFFF;
rommem[24225] <= 16'hFFFF;
rommem[24226] <= 16'hFFFF;
rommem[24227] <= 16'hFFFF;
rommem[24228] <= 16'hFFFF;
rommem[24229] <= 16'hFFFF;
rommem[24230] <= 16'hFFFF;
rommem[24231] <= 16'hFFFF;
rommem[24232] <= 16'hFFFF;
rommem[24233] <= 16'hFFFF;
rommem[24234] <= 16'hFFFF;
rommem[24235] <= 16'hFFFF;
rommem[24236] <= 16'hFFFF;
rommem[24237] <= 16'hFFFF;
rommem[24238] <= 16'hFFFF;
rommem[24239] <= 16'hFFFF;
rommem[24240] <= 16'hFFFF;
rommem[24241] <= 16'hFFFF;
rommem[24242] <= 16'hFFFF;
rommem[24243] <= 16'hFFFF;
rommem[24244] <= 16'hFFFF;
rommem[24245] <= 16'hFFFF;
rommem[24246] <= 16'hFFFF;
rommem[24247] <= 16'hFFFF;
rommem[24248] <= 16'hFFFF;
rommem[24249] <= 16'hFFFF;
rommem[24250] <= 16'hFFFF;
rommem[24251] <= 16'hFFFF;
rommem[24252] <= 16'hFFFF;
rommem[24253] <= 16'hFFFF;
rommem[24254] <= 16'hFFFF;
rommem[24255] <= 16'hFFFF;
rommem[24256] <= 16'hFFFF;
rommem[24257] <= 16'hFFFF;
rommem[24258] <= 16'hFFFF;
rommem[24259] <= 16'hFFFF;
rommem[24260] <= 16'hFFFF;
rommem[24261] <= 16'hFFFF;
rommem[24262] <= 16'hFFFF;
rommem[24263] <= 16'hFFFF;
rommem[24264] <= 16'hFFFF;
rommem[24265] <= 16'hFFFF;
rommem[24266] <= 16'hFFFF;
rommem[24267] <= 16'hFFFF;
rommem[24268] <= 16'hFFFF;
rommem[24269] <= 16'hFFFF;
rommem[24270] <= 16'hFFFF;
rommem[24271] <= 16'hFFFF;
rommem[24272] <= 16'hFFFF;
rommem[24273] <= 16'hFFFF;
rommem[24274] <= 16'hFFFF;
rommem[24275] <= 16'hFFFF;
rommem[24276] <= 16'hFFFF;
rommem[24277] <= 16'hFFFF;
rommem[24278] <= 16'hFFFF;
rommem[24279] <= 16'hFFFF;
rommem[24280] <= 16'hFFFF;
rommem[24281] <= 16'hFFFF;
rommem[24282] <= 16'hFFFF;
rommem[24283] <= 16'hFFFF;
rommem[24284] <= 16'hFFFF;
rommem[24285] <= 16'hFFFF;
rommem[24286] <= 16'hFFFF;
rommem[24287] <= 16'hFFFF;
rommem[24288] <= 16'hFFFF;
rommem[24289] <= 16'hFFFF;
rommem[24290] <= 16'hFFFF;
rommem[24291] <= 16'hFFFF;
rommem[24292] <= 16'hFFFF;
rommem[24293] <= 16'hFFFF;
rommem[24294] <= 16'hFFFF;
rommem[24295] <= 16'hFFFF;
rommem[24296] <= 16'hFFFF;
rommem[24297] <= 16'hFFFF;
rommem[24298] <= 16'hFFFF;
rommem[24299] <= 16'hFFFF;
rommem[24300] <= 16'hFFFF;
rommem[24301] <= 16'hFFFF;
rommem[24302] <= 16'hFFFF;
rommem[24303] <= 16'hFFFF;
rommem[24304] <= 16'hFFFF;
rommem[24305] <= 16'hFFFF;
rommem[24306] <= 16'hFFFF;
rommem[24307] <= 16'hFFFF;
rommem[24308] <= 16'hFFFF;
rommem[24309] <= 16'hFFFF;
rommem[24310] <= 16'hFFFF;
rommem[24311] <= 16'hFFFF;
rommem[24312] <= 16'hFFFF;
rommem[24313] <= 16'hFFFF;
rommem[24314] <= 16'hFFFF;
rommem[24315] <= 16'hFFFF;
rommem[24316] <= 16'hFFFF;
rommem[24317] <= 16'hFFFF;
rommem[24318] <= 16'hFFFF;
rommem[24319] <= 16'hFFFF;
rommem[24320] <= 16'hFFFF;
rommem[24321] <= 16'hFFFF;
rommem[24322] <= 16'hFFFF;
rommem[24323] <= 16'hFFFF;
rommem[24324] <= 16'hFFFF;
rommem[24325] <= 16'hFFFF;
rommem[24326] <= 16'hFFFF;
rommem[24327] <= 16'hFFFF;
rommem[24328] <= 16'hFFFF;
rommem[24329] <= 16'hFFFF;
rommem[24330] <= 16'hFFFF;
rommem[24331] <= 16'hFFFF;
rommem[24332] <= 16'hFFFF;
rommem[24333] <= 16'hFFFF;
rommem[24334] <= 16'hFFFF;
rommem[24335] <= 16'hFFFF;
rommem[24336] <= 16'hFFFF;
rommem[24337] <= 16'hFFFF;
rommem[24338] <= 16'hFFFF;
rommem[24339] <= 16'hFFFF;
rommem[24340] <= 16'hFFFF;
rommem[24341] <= 16'hFFFF;
rommem[24342] <= 16'hFFFF;
rommem[24343] <= 16'hFFFF;
rommem[24344] <= 16'hFFFF;
rommem[24345] <= 16'hFFFF;
rommem[24346] <= 16'hFFFF;
rommem[24347] <= 16'hFFFF;
rommem[24348] <= 16'hFFFF;
rommem[24349] <= 16'hFFFF;
rommem[24350] <= 16'hFFFF;
rommem[24351] <= 16'hFFFF;
rommem[24352] <= 16'hFFFF;
rommem[24353] <= 16'hFFFF;
rommem[24354] <= 16'hFFFF;
rommem[24355] <= 16'hFFFF;
rommem[24356] <= 16'hFFFF;
rommem[24357] <= 16'hFFFF;
rommem[24358] <= 16'hFFFF;
rommem[24359] <= 16'hFFFF;
rommem[24360] <= 16'hFFFF;
rommem[24361] <= 16'hFFFF;
rommem[24362] <= 16'hFFFF;
rommem[24363] <= 16'hFFFF;
rommem[24364] <= 16'hFFFF;
rommem[24365] <= 16'hFFFF;
rommem[24366] <= 16'hFFFF;
rommem[24367] <= 16'hFFFF;
rommem[24368] <= 16'hFFFF;
rommem[24369] <= 16'hFFFF;
rommem[24370] <= 16'hFFFF;
rommem[24371] <= 16'hFFFF;
rommem[24372] <= 16'hFFFF;
rommem[24373] <= 16'hFFFF;
rommem[24374] <= 16'hFFFF;
rommem[24375] <= 16'hFFFF;
rommem[24376] <= 16'hFFFF;
rommem[24377] <= 16'hFFFF;
rommem[24378] <= 16'hFFFF;
rommem[24379] <= 16'hFFFF;
rommem[24380] <= 16'hFFFF;
rommem[24381] <= 16'hFFFF;
rommem[24382] <= 16'hFFFF;
rommem[24383] <= 16'hFFFF;
rommem[24384] <= 16'hFFFF;
rommem[24385] <= 16'hFFFF;
rommem[24386] <= 16'hFFFF;
rommem[24387] <= 16'hFFFF;
rommem[24388] <= 16'hFFFF;
rommem[24389] <= 16'hFFFF;
rommem[24390] <= 16'hFFFF;
rommem[24391] <= 16'hFFFF;
rommem[24392] <= 16'hFFFF;
rommem[24393] <= 16'hFFFF;
rommem[24394] <= 16'hFFFF;
rommem[24395] <= 16'hFFFF;
rommem[24396] <= 16'hFFFF;
rommem[24397] <= 16'hFFFF;
rommem[24398] <= 16'hFFFF;
rommem[24399] <= 16'hFFFF;
rommem[24400] <= 16'hFFFF;
rommem[24401] <= 16'hFFFF;
rommem[24402] <= 16'hFFFF;
rommem[24403] <= 16'hFFFF;
rommem[24404] <= 16'hFFFF;
rommem[24405] <= 16'hFFFF;
rommem[24406] <= 16'hFFFF;
rommem[24407] <= 16'hFFFF;
rommem[24408] <= 16'hFFFF;
rommem[24409] <= 16'hFFFF;
rommem[24410] <= 16'hFFFF;
rommem[24411] <= 16'hFFFF;
rommem[24412] <= 16'hFFFF;
rommem[24413] <= 16'hFFFF;
rommem[24414] <= 16'hFFFF;
rommem[24415] <= 16'hFFFF;
rommem[24416] <= 16'hFFFF;
rommem[24417] <= 16'hFFFF;
rommem[24418] <= 16'hFFFF;
rommem[24419] <= 16'hFFFF;
rommem[24420] <= 16'hFFFF;
rommem[24421] <= 16'hFFFF;
rommem[24422] <= 16'hFFFF;
rommem[24423] <= 16'hFFFF;
rommem[24424] <= 16'hFFFF;
rommem[24425] <= 16'hFFFF;
rommem[24426] <= 16'hFFFF;
rommem[24427] <= 16'hFFFF;
rommem[24428] <= 16'hFFFF;
rommem[24429] <= 16'hFFFF;
rommem[24430] <= 16'hFFFF;
rommem[24431] <= 16'hFFFF;
rommem[24432] <= 16'hFFFF;
rommem[24433] <= 16'hFFFF;
rommem[24434] <= 16'hFFFF;
rommem[24435] <= 16'hFFFF;
rommem[24436] <= 16'hFFFF;
rommem[24437] <= 16'hFFFF;
rommem[24438] <= 16'hFFFF;
rommem[24439] <= 16'hFFFF;
rommem[24440] <= 16'hFFFF;
rommem[24441] <= 16'hFFFF;
rommem[24442] <= 16'hFFFF;
rommem[24443] <= 16'hFFFF;
rommem[24444] <= 16'hFFFF;
rommem[24445] <= 16'hFFFF;
rommem[24446] <= 16'hFFFF;
rommem[24447] <= 16'hFFFF;
rommem[24448] <= 16'hFFFF;
rommem[24449] <= 16'hFFFF;
rommem[24450] <= 16'hFFFF;
rommem[24451] <= 16'hFFFF;
rommem[24452] <= 16'hFFFF;
rommem[24453] <= 16'hFFFF;
rommem[24454] <= 16'hFFFF;
rommem[24455] <= 16'hFFFF;
rommem[24456] <= 16'hFFFF;
rommem[24457] <= 16'hFFFF;
rommem[24458] <= 16'hFFFF;
rommem[24459] <= 16'hFFFF;
rommem[24460] <= 16'hFFFF;
rommem[24461] <= 16'hFFFF;
rommem[24462] <= 16'hFFFF;
rommem[24463] <= 16'hFFFF;
rommem[24464] <= 16'hFFFF;
rommem[24465] <= 16'hFFFF;
rommem[24466] <= 16'hFFFF;
rommem[24467] <= 16'hFFFF;
rommem[24468] <= 16'hFFFF;
rommem[24469] <= 16'hFFFF;
rommem[24470] <= 16'hFFFF;
rommem[24471] <= 16'hFFFF;
rommem[24472] <= 16'hFFFF;
rommem[24473] <= 16'hFFFF;
rommem[24474] <= 16'hFFFF;
rommem[24475] <= 16'hFFFF;
rommem[24476] <= 16'hFFFF;
rommem[24477] <= 16'hFFFF;
rommem[24478] <= 16'hFFFF;
rommem[24479] <= 16'hFFFF;
rommem[24480] <= 16'hFFFF;
rommem[24481] <= 16'hFFFF;
rommem[24482] <= 16'hFFFF;
rommem[24483] <= 16'hFFFF;
rommem[24484] <= 16'hFFFF;
rommem[24485] <= 16'hFFFF;
rommem[24486] <= 16'hFFFF;
rommem[24487] <= 16'hFFFF;
rommem[24488] <= 16'hFFFF;
rommem[24489] <= 16'hFFFF;
rommem[24490] <= 16'hFFFF;
rommem[24491] <= 16'hFFFF;
rommem[24492] <= 16'hFFFF;
rommem[24493] <= 16'hFFFF;
rommem[24494] <= 16'hFFFF;
rommem[24495] <= 16'hFFFF;
rommem[24496] <= 16'hFFFF;
rommem[24497] <= 16'hFFFF;
rommem[24498] <= 16'hFFFF;
rommem[24499] <= 16'hFFFF;
rommem[24500] <= 16'hFFFF;
rommem[24501] <= 16'hFFFF;
rommem[24502] <= 16'hFFFF;
rommem[24503] <= 16'hFFFF;
rommem[24504] <= 16'hFFFF;
rommem[24505] <= 16'hFFFF;
rommem[24506] <= 16'hFFFF;
rommem[24507] <= 16'hFFFF;
rommem[24508] <= 16'hFFFF;
rommem[24509] <= 16'hFFFF;
rommem[24510] <= 16'hFFFF;
rommem[24511] <= 16'hFFFF;
rommem[24512] <= 16'hFFFF;
rommem[24513] <= 16'hFFFF;
rommem[24514] <= 16'hFFFF;
rommem[24515] <= 16'hFFFF;
rommem[24516] <= 16'hFFFF;
rommem[24517] <= 16'hFFFF;
rommem[24518] <= 16'hFFFF;
rommem[24519] <= 16'hFFFF;
rommem[24520] <= 16'hFFFF;
rommem[24521] <= 16'hFFFF;
rommem[24522] <= 16'hFFFF;
rommem[24523] <= 16'hFFFF;
rommem[24524] <= 16'hFFFF;
rommem[24525] <= 16'hFFFF;
rommem[24526] <= 16'hFFFF;
rommem[24527] <= 16'hFFFF;
rommem[24528] <= 16'hFFFF;
rommem[24529] <= 16'hFFFF;
rommem[24530] <= 16'hFFFF;
rommem[24531] <= 16'hFFFF;
rommem[24532] <= 16'hFFFF;
rommem[24533] <= 16'hFFFF;
rommem[24534] <= 16'hFFFF;
rommem[24535] <= 16'hFFFF;
rommem[24536] <= 16'hFFFF;
rommem[24537] <= 16'hFFFF;
rommem[24538] <= 16'hFFFF;
rommem[24539] <= 16'hFFFF;
rommem[24540] <= 16'hFFFF;
rommem[24541] <= 16'hFFFF;
rommem[24542] <= 16'hFFFF;
rommem[24543] <= 16'hFFFF;
rommem[24544] <= 16'hFFFF;
rommem[24545] <= 16'hFFFF;
rommem[24546] <= 16'hFFFF;
rommem[24547] <= 16'hFFFF;
rommem[24548] <= 16'hFFFF;
rommem[24549] <= 16'hFFFF;
rommem[24550] <= 16'hFFFF;
rommem[24551] <= 16'hFFFF;
rommem[24552] <= 16'hFFFF;
rommem[24553] <= 16'hFFFF;
rommem[24554] <= 16'hFFFF;
rommem[24555] <= 16'hFFFF;
rommem[24556] <= 16'hFFFF;
rommem[24557] <= 16'hFFFF;
rommem[24558] <= 16'hFFFF;
rommem[24559] <= 16'hFFFF;
rommem[24560] <= 16'hFFFF;
rommem[24561] <= 16'hFFFF;
rommem[24562] <= 16'hFFFF;
rommem[24563] <= 16'hFFFF;
rommem[24564] <= 16'hFFFF;
rommem[24565] <= 16'hFFFF;
rommem[24566] <= 16'hFFFF;
rommem[24567] <= 16'hFFFF;
rommem[24568] <= 16'hFFFF;
rommem[24569] <= 16'hFFFF;
rommem[24570] <= 16'hFFFF;
rommem[24571] <= 16'hFFFF;
rommem[24572] <= 16'hFFFF;
rommem[24573] <= 16'hFFFF;
rommem[24574] <= 16'hFFFF;
rommem[24575] <= 16'hFFFF;
rommem[24576] <= 16'h6000;
rommem[24577] <= 16'h0022;
rommem[24578] <= 16'h6000;
rommem[24579] <= 16'h005A;
rommem[24580] <= 16'h6000;
rommem[24581] <= 16'h0B68;
rommem[24582] <= 16'h6000;
rommem[24583] <= 16'h0B74;
rommem[24584] <= 16'h6000;
rommem[24585] <= 16'h0B86;
rommem[24586] <= 16'h6000;
rommem[24587] <= 16'h0B94;
rommem[24588] <= 16'h6000;
rommem[24589] <= 16'h0BA6;
rommem[24590] <= 16'h0020;
rommem[24591] <= 16'h0000;
rommem[24592] <= 16'h1F00;
rommem[24593] <= 16'h0000;
rommem[24594] <= 16'h41F9;
rommem[24595] <= 16'hFFFC;
rommem[24596] <= 16'hC000;
rommem[24597] <= 16'h21C8;
rommem[24598] <= 16'h0600;
rommem[24599] <= 16'h2E79;
rommem[24600] <= 16'hFFFC;
rommem[24601] <= 16'hC020;
rommem[24602] <= 16'h4DF9;
rommem[24603] <= 16'hFFFC;
rommem[24604] <= 16'hCBC6;
rommem[24605] <= 16'h6100;
rommem[24606] <= 16'h0B2A;
rommem[24607] <= 16'h21F9;
rommem[24608] <= 16'hFFFC;
rommem[24609] <= 16'hC01C;
rommem[24610] <= 16'h0624;
rommem[24611] <= 16'h2039;
rommem[24612] <= 16'hFFFC;
rommem[24613] <= 16'hC020;
rommem[24614] <= 16'h0480;
rommem[24615] <= 16'h0000;
rommem[24616] <= 16'h0800;
rommem[24617] <= 16'h21C0;
rommem[24618] <= 16'h062C;
rommem[24619] <= 16'h0480;
rommem[24620] <= 16'h0000;
rommem[24621] <= 16'h006C;
rommem[24622] <= 16'h21C0;
rommem[24623] <= 16'h0628;
rommem[24624] <= 16'h4280;
rommem[24625] <= 16'h21C0;
rommem[24626] <= 16'h0610;
rommem[24627] <= 16'h21C0;
rommem[24628] <= 16'h0608;
rommem[24629] <= 16'h21C0;
rommem[24630] <= 16'h0604;
rommem[24631] <= 16'h2E79;
rommem[24632] <= 16'hFFFC;
rommem[24633] <= 16'hC020;
rommem[24634] <= 16'h4DF9;
rommem[24635] <= 16'hFFFC;
rommem[24636] <= 16'hCBD1;
rommem[24637] <= 16'h6100;
rommem[24638] <= 16'h0AEA;
rommem[24639] <= 16'h103C;
rommem[24640] <= 16'h003E;
rommem[24641] <= 16'h6100;
rommem[24642] <= 16'h0810;
rommem[24643] <= 16'h6100;
rommem[24644] <= 16'h0A7A;
rommem[24645] <= 16'h2848;
rommem[24646] <= 16'h41F8;
rommem[24647] <= 16'h0630;
rommem[24648] <= 16'h6100;
rommem[24649] <= 16'h0A2C;
rommem[24650] <= 16'h6100;
rommem[24651] <= 16'h0A60;
rommem[24652] <= 16'h4A81;
rommem[24653] <= 16'h6700;
rommem[24654] <= 16'h011A;
rommem[24655] <= 16'hB2BC;
rommem[24656] <= 16'h0000;
rommem[24657] <= 16'hFFFF;
rommem[24658] <= 16'h6400;
rommem[24659] <= 16'h07E4;
rommem[24660] <= 16'h1101;
rommem[24661] <= 16'hE099;
rommem[24662] <= 16'h1101;
rommem[24663] <= 16'hE199;
rommem[24664] <= 16'h6100;
rommem[24665] <= 16'h0882;
rommem[24666] <= 16'h2A49;
rommem[24667] <= 16'h6612;
rommem[24668] <= 16'h6100;
rommem[24669] <= 16'h08A2;
rommem[24670] <= 16'h244D;
rommem[24671] <= 16'h2678;
rommem[24672] <= 16'h0624;
rommem[24673] <= 16'h6100;
rommem[24674] <= 16'h08A2;
rommem[24675] <= 16'h21CA;
rommem[24676] <= 16'h0624;
rommem[24677] <= 16'h200C;
rommem[24678] <= 16'h9088;
rommem[24679] <= 16'hB0BC;
rommem[24680] <= 16'h0000;
rommem[24681] <= 16'h0003;
rommem[24682] <= 16'h67A8;
rommem[24683] <= 16'h2678;
rommem[24684] <= 16'h0624;
rommem[24685] <= 16'h2C4B;
rommem[24686] <= 16'hD7C0;
rommem[24687] <= 16'h2038;
rommem[24688] <= 16'h0628;
rommem[24689] <= 16'hB08B;
rommem[24690] <= 16'h6300;
rommem[24691] <= 16'h079A;
rommem[24692] <= 16'h21CB;
rommem[24693] <= 16'h0624;
rommem[24694] <= 16'h224E;
rommem[24695] <= 16'h244D;
rommem[24696] <= 16'h6100;
rommem[24697] <= 16'h087E;
rommem[24698] <= 16'h2248;
rommem[24699] <= 16'h244D;
rommem[24700] <= 16'h264C;
rommem[24701] <= 16'h6100;
rommem[24702] <= 16'h086A;
rommem[24703] <= 16'h6000;
rommem[24704] <= 16'hFF7E;
rommem[24705] <= 16'h4C49;
rommem[24706] <= 16'h53D4;
rommem[24707] <= 16'h4C4F;
rommem[24708] <= 16'h41C4;
rommem[24709] <= 16'h4E45;
rommem[24710] <= 16'hD752;
rommem[24711] <= 16'h55CE;
rommem[24712] <= 16'h5341;
rommem[24713] <= 16'h56C5;
rommem[24714] <= 16'h4E45;
rommem[24715] <= 16'h58D4;
rommem[24716] <= 16'h4C45;
rommem[24717] <= 16'hD449;
rommem[24718] <= 16'hC647;
rommem[24719] <= 16'h4F54;
rommem[24720] <= 16'hCF47;
rommem[24721] <= 16'h4F53;
rommem[24722] <= 16'h55C2;
rommem[24723] <= 16'h5245;
rommem[24724] <= 16'h5455;
rommem[24725] <= 16'h52CE;
rommem[24726] <= 16'h5245;
rommem[24727] <= 16'hCD46;
rommem[24728] <= 16'h4FD2;
rommem[24729] <= 16'h494E;
rommem[24730] <= 16'h5055;
rommem[24731] <= 16'hD450;
rommem[24732] <= 16'h5249;
rommem[24733] <= 16'h4ED4;
rommem[24734] <= 16'h504F;
rommem[24735] <= 16'h4BC5;
rommem[24736] <= 16'h5354;
rommem[24737] <= 16'h4FD0;
rommem[24738] <= 16'h4259;
rommem[24739] <= 16'hC543;
rommem[24740] <= 16'h414C;
rommem[24741] <= 16'hCC00;
rommem[24742] <= 16'h5045;
rommem[24743] <= 16'h45CB;
rommem[24744] <= 16'h524E;
rommem[24745] <= 16'hC441;
rommem[24746] <= 16'h42D3;
rommem[24747] <= 16'h5349;
rommem[24748] <= 16'h5AC5;
rommem[24749] <= 16'h0054;
rommem[24750] <= 16'hCF00;
rommem[24751] <= 16'h5354;
rommem[24752] <= 16'h45D0;
rommem[24753] <= 16'h003E;
rommem[24754] <= 16'hBD3C;
rommem[24755] <= 16'hBEBE;
rommem[24756] <= 16'hBD3C;
rommem[24757] <= 16'hBDBC;
rommem[24758] <= 16'h0000;
rommem[24759] <= 16'hC266;
rommem[24760] <= 16'hC4A8;
rommem[24761] <= 16'hC200;
rommem[24762] <= 16'hC214;
rommem[24763] <= 16'hC50C;
rommem[24764] <= 16'hC3B4;
rommem[24765] <= 16'hC498;
rommem[24766] <= 16'hC404;
rommem[24767] <= 16'hC252;
rommem[24768] <= 16'hC2FC;
rommem[24769] <= 16'hC324;
rommem[24770] <= 16'hC402;
rommem[24771] <= 16'hC342;
rommem[24772] <= 16'hC42A;
rommem[24773] <= 16'hC292;
rommem[24774] <= 16'hC590;
rommem[24775] <= 16'hC20C;
rommem[24776] <= 16'hC018;
rommem[24777] <= 16'hC5AC;
rommem[24778] <= 16'hC492;
rommem[24779] <= 16'hC7A2;
rommem[24780] <= 16'hC7AE;
rommem[24781] <= 16'hC7E4;
rommem[24782] <= 16'hC7F4;
rommem[24783] <= 16'hC6A6;
rommem[24784] <= 16'hC35E;
rommem[24785] <= 16'hC83E;
rommem[24786] <= 16'hC376;
rommem[24787] <= 16'hC37C;
rommem[24788] <= 16'hC5D8;
rommem[24789] <= 16'hC5E0;
rommem[24790] <= 16'hC5E8;
rommem[24791] <= 16'hC5F8;
rommem[24792] <= 16'hC5F0;
rommem[24793] <= 16'hC602;
rommem[24794] <= 16'hC614;
rommem[24795] <= 16'h43F9;
rommem[24796] <= 16'hFFFC;
rommem[24797] <= 16'hC102;
rommem[24798] <= 16'h45F9;
rommem[24799] <= 16'hFFFC;
rommem[24800] <= 16'hC16E;
rommem[24801] <= 16'h6100;
rommem[24802] <= 16'h0932;
rommem[24803] <= 16'h2648;
rommem[24804] <= 16'h4202;
rommem[24805] <= 16'h1018;
rommem[24806] <= 16'h1211;
rommem[24807] <= 16'h6604;
rommem[24808] <= 16'h204B;
rommem[24809] <= 16'h6024;
rommem[24810] <= 16'h1600;
rommem[24811] <= 16'hC602;
rommem[24812] <= 16'hB63C;
rommem[24813] <= 16'h002E;
rommem[24814] <= 16'h671A;
rommem[24815] <= 16'h0201;
rommem[24816] <= 16'h007F;
rommem[24817] <= 16'hB200;
rommem[24818] <= 16'h670C;
rommem[24819] <= 16'h548A;
rommem[24820] <= 16'h204B;
rommem[24821] <= 16'h4202;
rommem[24822] <= 16'h4A19;
rommem[24823] <= 16'h6AFC;
rommem[24824] <= 16'h60D8;
rommem[24825] <= 16'h74FF;
rommem[24826] <= 16'h4A19;
rommem[24827] <= 16'h6AD2;
rommem[24828] <= 16'h47F8;
rommem[24829] <= 16'h0000;
rommem[24830] <= 16'h2652;
rommem[24831] <= 16'h4ED3;
rommem[24832] <= 16'h6100;
rommem[24833] <= 16'h0630;
rommem[24834] <= 16'h21F9;
rommem[24835] <= 16'hFFFC;
rommem[24836] <= 16'hC01C;
rommem[24837] <= 16'h0624;
rommem[24838] <= 16'h6100;
rommem[24839] <= 16'h0624;
rommem[24840] <= 16'h6000;
rommem[24841] <= 16'hFE4E;
rommem[24842] <= 16'h6100;
rommem[24843] <= 16'h061C;
rommem[24844] <= 16'h2079;
rommem[24845] <= 16'hFFFC;
rommem[24846] <= 16'hC01C;
rommem[24847] <= 16'h21C8;
rommem[24848] <= 16'h0604;
rommem[24849] <= 16'h4AB8;
rommem[24850] <= 16'h0604;
rommem[24851] <= 16'h6700;
rommem[24852] <= 16'hFE38;
rommem[24853] <= 16'h4281;
rommem[24854] <= 16'h2248;
rommem[24855] <= 16'h6100;
rommem[24856] <= 16'h0714;
rommem[24857] <= 16'h6500;
rommem[24858] <= 16'hFE2C;
rommem[24859] <= 16'h21C9;
rommem[24860] <= 16'h0604;
rommem[24861] <= 16'h2049;
rommem[24862] <= 16'h5488;
rommem[24863] <= 16'h6100;
rommem[24864] <= 16'h090E;
rommem[24865] <= 16'h43F9;
rommem[24866] <= 16'hFFFC;
rommem[24867] <= 16'hC114;
rommem[24868] <= 16'h45F9;
rommem[24869] <= 16'hFFFC;
rommem[24870] <= 16'hC178;
rommem[24871] <= 16'h6000;
rommem[24872] <= 16'hFF72;
rommem[24873] <= 16'h6100;
rommem[24874] <= 16'h036E;
rommem[24875] <= 16'h6100;
rommem[24876] <= 16'h05DA;
rommem[24877] <= 16'h2200;
rommem[24878] <= 16'h6100;
rommem[24879] <= 16'h06D6;
rommem[24880] <= 16'h6600;
rommem[24881] <= 16'h0628;
rommem[24882] <= 16'h60D0;
rommem[24883] <= 16'h6100;
rommem[24884] <= 16'h0856;
rommem[24885] <= 16'h6100;
rommem[24886] <= 16'h05C6;
rommem[24887] <= 16'h6100;
rommem[24888] <= 16'h06C4;
rommem[24889] <= 16'h6500;
rommem[24890] <= 16'hFDEC;
rommem[24891] <= 16'h6100;
rommem[24892] <= 16'h0810;
rommem[24893] <= 16'h6100;
rommem[24894] <= 16'h08D2;
rommem[24895] <= 16'h670C;
rommem[24896] <= 16'hB03C;
rommem[24897] <= 16'h0013;
rommem[24898] <= 16'h6606;
rommem[24899] <= 16'h6100;
rommem[24900] <= 16'h08C6;
rommem[24901] <= 16'h67FA;
rommem[24902] <= 16'h6100;
rommem[24903] <= 16'h06B6;
rommem[24904] <= 16'h60E0;
rommem[24905] <= 16'h780B;
rommem[24906] <= 16'h6100;
rommem[24907] <= 16'h080E;
rommem[24908] <= 16'h3A07;
rommem[24909] <= 16'h6100;
rommem[24910] <= 16'h08C4;
rommem[24911] <= 16'h609E;
rommem[24912] <= 16'h6100;
rommem[24913] <= 16'h0802;
rommem[24914] <= 16'h0D09;
rommem[24915] <= 16'h6100;
rommem[24916] <= 16'h08B8;
rommem[24917] <= 16'h6000;
rommem[24918] <= 16'hFF76;
rommem[24919] <= 16'h6100;
rommem[24920] <= 16'h07F4;
rommem[24921] <= 16'h2309;
rommem[24922] <= 16'h6100;
rommem[24923] <= 16'h030C;
rommem[24924] <= 16'h2800;
rommem[24925] <= 16'h6016;
rommem[24926] <= 16'h6100;
rommem[24927] <= 16'h07E6;
rommem[24928] <= 16'h240B;
rommem[24929] <= 16'h6100;
rommem[24930] <= 16'h02FE;
rommem[24931] <= 16'h6100;
rommem[24932] <= 16'hFD40;
rommem[24933] <= 16'h6006;
rommem[24934] <= 16'h6100;
rommem[24935] <= 16'h0706;
rommem[24936] <= 16'h6012;
rommem[24937] <= 16'h6100;
rommem[24938] <= 16'h07D0;
rommem[24939] <= 16'h2C07;
rommem[24940] <= 16'h6100;
rommem[24941] <= 16'h053E;
rommem[24942] <= 16'h60D0;
rommem[24943] <= 16'h6100;
rommem[24944] <= 16'h0880;
rommem[24945] <= 16'h6010;
rommem[24946] <= 16'h2F04;
rommem[24947] <= 16'h6100;
rommem[24948] <= 16'h02DA;
rommem[24949] <= 16'h281F;
rommem[24950] <= 16'h2200;
rommem[24951] <= 16'h6100;
rommem[24952] <= 16'h0724;
rommem[24953] <= 16'h60DE;
rommem[24954] <= 16'h6100;
rommem[24955] <= 16'h0522;
rommem[24956] <= 16'h6000;
rommem[24957] <= 16'h0544;
rommem[24958] <= 16'h6100;
rommem[24959] <= 16'h0694;
rommem[24960] <= 16'h6100;
rommem[24961] <= 16'h02C0;
rommem[24962] <= 16'h2F08;
rommem[24963] <= 16'h2200;
rommem[24964] <= 16'h6100;
rommem[24965] <= 16'h062A;
rommem[24966] <= 16'h6600;
rommem[24967] <= 16'h057E;
rommem[24968] <= 16'h2F38;
rommem[24969] <= 16'h0604;
rommem[24970] <= 16'h2F38;
rommem[24971] <= 16'h0608;
rommem[24972] <= 16'h42B8;
rommem[24973] <= 16'h0610;
rommem[24974] <= 16'h21CF;
rommem[24975] <= 16'h0608;
rommem[24976] <= 16'h6000;
rommem[24977] <= 16'hFF14;
rommem[24978] <= 16'h6100;
rommem[24979] <= 16'h050C;
rommem[24980] <= 16'h2238;
rommem[24981] <= 16'h0608;
rommem[24982] <= 16'h6700;
rommem[24983] <= 16'h0510;
rommem[24984] <= 16'h2E41;
rommem[24985] <= 16'h21DF;
rommem[24986] <= 16'h0608;
rommem[24987] <= 16'h21DF;
rommem[24988] <= 16'h0604;
rommem[24989] <= 16'h205F;
rommem[24990] <= 16'h6100;
rommem[24991] <= 16'h063A;
rommem[24992] <= 16'h60B2;
rommem[24993] <= 16'h6100;
rommem[24994] <= 16'h064E;
rommem[24995] <= 16'h6100;
rommem[24996] <= 16'h04B6;
rommem[24997] <= 16'h21CE;
rommem[24998] <= 16'h0610;
rommem[24999] <= 16'h43F9;
rommem[25000] <= 16'hFFFC;
rommem[25001] <= 16'hC15B;
rommem[25002] <= 16'h45F9;
rommem[25003] <= 16'hFFFC;
rommem[25004] <= 16'hC1A0;
rommem[25005] <= 16'h6000;
rommem[25006] <= 16'hFE66;
rommem[25007] <= 16'h6100;
rommem[25008] <= 16'h0262;
rommem[25009] <= 16'h21C0;
rommem[25010] <= 16'h0618;
rommem[25011] <= 16'h43F9;
rommem[25012] <= 16'hFFFC;
rommem[25013] <= 16'hC15E;
rommem[25014] <= 16'h45F9;
rommem[25015] <= 16'hFFFC;
rommem[25016] <= 16'hC1A4;
rommem[25017] <= 16'h6000;
rommem[25018] <= 16'hFE4E;
rommem[25019] <= 16'h6100;
rommem[25020] <= 16'h024A;
rommem[25021] <= 16'h6002;
rommem[25022] <= 16'h7001;
rommem[25023] <= 16'h21C0;
rommem[25024] <= 16'h0614;
rommem[25025] <= 16'h21F8;
rommem[25026] <= 16'h0604;
rommem[25027] <= 16'h061C;
rommem[25028] <= 16'h21C8;
rommem[25029] <= 16'h0620;
rommem[25030] <= 16'h2C4F;
rommem[25031] <= 16'h6006;
rommem[25032] <= 16'hDDFC;
rommem[25033] <= 16'h0000;
rommem[25034] <= 16'h0014;
rommem[25035] <= 16'h2016;
rommem[25036] <= 16'h6716;
rommem[25037] <= 16'hB0B8;
rommem[25038] <= 16'h0610;
rommem[25039] <= 16'h66F0;
rommem[25040] <= 16'h244F;
rommem[25041] <= 16'h224E;
rommem[25042] <= 16'h47F8;
rommem[25043] <= 16'h0014;
rommem[25044] <= 16'hD7C9;
rommem[25045] <= 16'h6100;
rommem[25046] <= 16'h05C4;
rommem[25047] <= 16'h2E4B;
rommem[25048] <= 16'h6000;
rommem[25049] <= 16'hFF42;
rommem[25050] <= 16'h6100;
rommem[25051] <= 16'h031E;
rommem[25052] <= 16'h6500;
rommem[25053] <= 16'h0484;
rommem[25054] <= 16'h2240;
rommem[25055] <= 16'h2038;
rommem[25056] <= 16'h0610;
rommem[25057] <= 16'h6700;
rommem[25058] <= 16'h047A;
rommem[25059] <= 16'hB3C0;
rommem[25060] <= 16'h6706;
rommem[25061] <= 16'h6100;
rommem[25062] <= 16'h05AC;
rommem[25063] <= 16'h60EE;
rommem[25064] <= 16'h2011;
rommem[25065] <= 16'hD0B8;
rommem[25066] <= 16'h0614;
rommem[25067] <= 16'h6900;
rommem[25068] <= 16'h04B2;
rommem[25069] <= 16'h2280;
rommem[25070] <= 16'h2238;
rommem[25071] <= 16'h0618;
rommem[25072] <= 16'h4AB8;
rommem[25073] <= 16'h0614;
rommem[25074] <= 16'h6A02;
rommem[25075] <= 16'hC141;
rommem[25076] <= 16'hB280;
rommem[25077] <= 16'h6D0E;
rommem[25078] <= 16'h21F8;
rommem[25079] <= 16'h061C;
rommem[25080] <= 16'h0604;
rommem[25081] <= 16'h2078;
rommem[25082] <= 16'h0620;
rommem[25083] <= 16'h6000;
rommem[25084] <= 16'hFEFC;
rommem[25085] <= 16'h6100;
rommem[25086] <= 16'h057C;
rommem[25087] <= 16'h6000;
rommem[25088] <= 16'hFEF4;
rommem[25089] <= 16'h600A;
rommem[25090] <= 16'h6100;
rommem[25091] <= 16'h01BC;
rommem[25092] <= 16'h4A80;
rommem[25093] <= 16'h6600;
rommem[25094] <= 16'hFE32;
rommem[25095] <= 16'h2248;
rommem[25096] <= 16'h4281;
rommem[25097] <= 16'h6100;
rommem[25098] <= 16'h054A;
rommem[25099] <= 16'h6400;
rommem[25100] <= 16'hFE1E;
rommem[25101] <= 16'h6000;
rommem[25102] <= 16'hFC44;
rommem[25103] <= 16'h2E78;
rommem[25104] <= 16'h060C;
rommem[25105] <= 16'h21DF;
rommem[25106] <= 16'h0604;
rommem[25107] <= 16'h588F;
rommem[25108] <= 16'h205F;
rommem[25109] <= 16'h2F08;
rommem[25110] <= 16'h6100;
rommem[25111] <= 16'h05A6;
rommem[25112] <= 16'h600A;
rommem[25113] <= 16'h6100;
rommem[25114] <= 16'h02A0;
rommem[25115] <= 16'h654C;
rommem[25116] <= 16'h2440;
rommem[25117] <= 16'h601A;
rommem[25118] <= 16'h2F08;
rommem[25119] <= 16'h6100;
rommem[25120] <= 16'h0294;
rommem[25121] <= 16'h6500;
rommem[25122] <= 16'h03FA;
rommem[25123] <= 16'h2440;
rommem[25124] <= 16'h1410;
rommem[25125] <= 16'h4200;
rommem[25126] <= 16'h1080;
rommem[25127] <= 16'h225F;
rommem[25128] <= 16'h6100;
rommem[25129] <= 16'h0566;
rommem[25130] <= 16'h1082;
rommem[25131] <= 16'h2F08;
rommem[25132] <= 16'h2F38;
rommem[25133] <= 16'h0604;
rommem[25134] <= 16'h21FC;
rommem[25135] <= 16'hFFFF;
rommem[25136] <= 16'hFFFF;
rommem[25137] <= 16'h0604;
rommem[25138] <= 16'h21CF;
rommem[25139] <= 16'h060C;
rommem[25140] <= 16'h2F0A;
rommem[25141] <= 16'h103C;
rommem[25142] <= 16'h003A;
rommem[25143] <= 16'h6100;
rommem[25144] <= 16'h0424;
rommem[25145] <= 16'h41F8;
rommem[25146] <= 16'h0630;
rommem[25147] <= 16'h6100;
rommem[25148] <= 16'h014A;
rommem[25149] <= 16'h245F;
rommem[25150] <= 16'h2480;
rommem[25151] <= 16'h21DF;
rommem[25152] <= 16'h0604;
rommem[25153] <= 16'h205F;
rommem[25154] <= 16'h588F;
rommem[25155] <= 16'h6100;
rommem[25156] <= 16'h061C;
rommem[25157] <= 16'h2C03;
rommem[25158] <= 16'h609C;
rommem[25159] <= 16'h6000;
rommem[25160] <= 16'hFE64;
rommem[25161] <= 16'h0C10;
rommem[25162] <= 16'h000D;
rommem[25163] <= 16'h670C;
rommem[25164] <= 16'h6100;
rommem[25165] <= 16'h0364;
rommem[25166] <= 16'h6100;
rommem[25167] <= 16'h0606;
rommem[25168] <= 16'h2C03;
rommem[25169] <= 16'h60F4;
rommem[25170] <= 16'h6000;
rommem[25171] <= 16'hFE4E;
rommem[25172] <= 16'h2079;
rommem[25173] <= 16'hFFFC;
rommem[25174] <= 16'hC01C;
rommem[25175] <= 16'h103C;
rommem[25176] <= 16'h000D;
rommem[25177] <= 16'h6100;
rommem[25178] <= 16'hFB5C;
rommem[25179] <= 16'h6100;
rommem[25180] <= 16'hFB5C;
rommem[25181] <= 16'h67FA;
rommem[25182] <= 16'hB03C;
rommem[25183] <= 16'h0040;
rommem[25184] <= 16'h6722;
rommem[25185] <= 16'hB03C;
rommem[25186] <= 16'h003A;
rommem[25187] <= 16'h66EE;
rommem[25188] <= 16'h6100;
rommem[25189] <= 16'h0022;
rommem[25190] <= 16'h10C1;
rommem[25191] <= 16'h6100;
rommem[25192] <= 16'h001C;
rommem[25193] <= 16'h10C1;
rommem[25194] <= 16'h6100;
rommem[25195] <= 16'hFB3E;
rommem[25196] <= 16'h67FA;
rommem[25197] <= 16'h10C0;
rommem[25198] <= 16'hB03C;
rommem[25199] <= 16'h000D;
rommem[25200] <= 16'h66F2;
rommem[25201] <= 16'h60D2;
rommem[25202] <= 16'h21C8;
rommem[25203] <= 16'h0624;
rommem[25204] <= 16'h6000;
rommem[25205] <= 16'hFB76;
rommem[25206] <= 16'h7401;
rommem[25207] <= 16'h4281;
rommem[25208] <= 16'h6100;
rommem[25209] <= 16'hFB22;
rommem[25210] <= 16'h67FA;
rommem[25211] <= 16'hB03C;
rommem[25212] <= 16'h0041;
rommem[25213] <= 16'h6502;
rommem[25214] <= 16'h5F00;
rommem[25215] <= 16'h0200;
rommem[25216] <= 16'h000F;
rommem[25217] <= 16'hE909;
rommem[25218] <= 16'h8200;
rommem[25219] <= 16'h51CA;
rommem[25220] <= 16'hFFE8;
rommem[25221] <= 16'h4E75;
rommem[25222] <= 16'h2079;
rommem[25223] <= 16'hFFFC;
rommem[25224] <= 16'hC01C;
rommem[25225] <= 16'h2278;
rommem[25226] <= 16'h0624;
rommem[25227] <= 16'h103C;
rommem[25228] <= 16'h000D;
rommem[25229] <= 16'h6100;
rommem[25230] <= 16'hFAF4;
rommem[25231] <= 16'h103C;
rommem[25232] <= 16'h000A;
rommem[25233] <= 16'h6100;
rommem[25234] <= 16'hFAEC;
rommem[25235] <= 16'hB3C8;
rommem[25236] <= 16'h6322;
rommem[25237] <= 16'h103C;
rommem[25238] <= 16'h003A;
rommem[25239] <= 16'h6100;
rommem[25240] <= 16'hFAE0;
rommem[25241] <= 16'h1218;
rommem[25242] <= 16'h6100;
rommem[25243] <= 16'h003A;
rommem[25244] <= 16'h1218;
rommem[25245] <= 16'h6100;
rommem[25246] <= 16'h0034;
rommem[25247] <= 16'h1018;
rommem[25248] <= 16'hB03C;
rommem[25249] <= 16'h000D;
rommem[25250] <= 16'h67D0;
rommem[25251] <= 16'h6100;
rommem[25252] <= 16'hFAC8;
rommem[25253] <= 16'h60F2;
rommem[25254] <= 16'h103C;
rommem[25255] <= 16'h0040;
rommem[25256] <= 16'h6100;
rommem[25257] <= 16'hFABE;
rommem[25258] <= 16'h103C;
rommem[25259] <= 16'h000D;
rommem[25260] <= 16'h6100;
rommem[25261] <= 16'hFAB6;
rommem[25262] <= 16'h103C;
rommem[25263] <= 16'h000A;
rommem[25264] <= 16'h6100;
rommem[25265] <= 16'hFAAE;
rommem[25266] <= 16'h103C;
rommem[25267] <= 16'h001A;
rommem[25268] <= 16'h6100;
rommem[25269] <= 16'hFAA6;
rommem[25270] <= 16'h6000;
rommem[25271] <= 16'hFAF2;
rommem[25272] <= 16'h7401;
rommem[25273] <= 16'hE919;
rommem[25274] <= 16'h1001;
rommem[25275] <= 16'h0200;
rommem[25276] <= 16'h000F;
rommem[25277] <= 16'h0600;
rommem[25278] <= 16'h0030;
rommem[25279] <= 16'hB03C;
rommem[25280] <= 16'h0039;
rommem[25281] <= 16'h6302;
rommem[25282] <= 16'h5E00;
rommem[25283] <= 16'h6100;
rommem[25284] <= 16'hFA88;
rommem[25285] <= 16'h51CA;
rommem[25286] <= 16'hFFE6;
rommem[25287] <= 16'h4E75;
rommem[25288] <= 16'h6100;
rommem[25289] <= 16'h0030;
rommem[25290] <= 16'h6100;
rommem[25291] <= 16'h050E;
rommem[25292] <= 16'h2C0F;
rommem[25293] <= 16'h2F00;
rommem[25294] <= 16'h6100;
rommem[25295] <= 16'h0024;
rommem[25296] <= 16'h225F;
rommem[25297] <= 16'h1280;
rommem[25298] <= 16'h6000;
rommem[25299] <= 16'hFD4E;
rommem[25300] <= 16'h6000;
rommem[25301] <= 16'h0294;
rommem[25302] <= 16'h6100;
rommem[25303] <= 16'h0014;
rommem[25304] <= 16'h4A80;
rommem[25305] <= 16'h6700;
rommem[25306] <= 16'h02D6;
rommem[25307] <= 16'h2F08;
rommem[25308] <= 16'h2240;
rommem[25309] <= 16'h4E91;
rommem[25310] <= 16'h205F;
rommem[25311] <= 16'h6000;
rommem[25312] <= 16'hFD34;
rommem[25313] <= 16'h6100;
rommem[25314] <= 16'h0066;
rommem[25315] <= 16'h2F00;
rommem[25316] <= 16'h43F9;
rommem[25317] <= 16'hFFFC;
rommem[25318] <= 16'hC163;
rommem[25319] <= 16'h45F9;
rommem[25320] <= 16'hFFFC;
rommem[25321] <= 16'hC1A8;
rommem[25322] <= 16'h6000;
rommem[25323] <= 16'hFBEC;
rommem[25324] <= 16'h6100;
rommem[25325] <= 16'h003E;
rommem[25326] <= 16'h6D2E;
rommem[25327] <= 16'h6030;
rommem[25328] <= 16'h6100;
rommem[25329] <= 16'h0036;
rommem[25330] <= 16'h6726;
rommem[25331] <= 16'h6028;
rommem[25332] <= 16'h6100;
rommem[25333] <= 16'h002E;
rommem[25334] <= 16'h6F1E;
rommem[25335] <= 16'h6020;
rommem[25336] <= 16'h6100;
rommem[25337] <= 16'h0026;
rommem[25338] <= 16'h6E16;
rommem[25339] <= 16'h6018;
rommem[25340] <= 16'h6100;
rommem[25341] <= 16'h001E;
rommem[25342] <= 16'h660E;
rommem[25343] <= 16'h6010;
rommem[25344] <= 16'h4E75;
rommem[25345] <= 16'h6100;
rommem[25346] <= 16'h0014;
rommem[25347] <= 16'h6C04;
rommem[25348] <= 16'h6006;
rommem[25349] <= 16'h4E75;
rommem[25350] <= 16'h4280;
rommem[25351] <= 16'h4E75;
rommem[25352] <= 16'h7001;
rommem[25353] <= 16'h4E75;
rommem[25354] <= 16'h201F;
rommem[25355] <= 16'h4E75;
rommem[25356] <= 16'h201F;
rommem[25357] <= 16'h221F;
rommem[25358] <= 16'h2F00;
rommem[25359] <= 16'h2F01;
rommem[25360] <= 16'h6100;
rommem[25361] <= 16'h0008;
rommem[25362] <= 16'h221F;
rommem[25363] <= 16'hB280;
rommem[25364] <= 16'h4E75;
rommem[25365] <= 16'h6100;
rommem[25366] <= 16'h0478;
rommem[25367] <= 16'h2D05;
rommem[25368] <= 16'h4280;
rommem[25369] <= 16'h6026;
rommem[25370] <= 16'h6100;
rommem[25371] <= 16'h046E;
rommem[25372] <= 16'h2B01;
rommem[25373] <= 16'h6100;
rommem[25374] <= 16'h002C;
rommem[25375] <= 16'h6100;
rommem[25376] <= 16'h0464;
rommem[25377] <= 16'h2B11;
rommem[25378] <= 16'h2F00;
rommem[25379] <= 16'h6100;
rommem[25380] <= 16'h0020;
rommem[25381] <= 16'h221F;
rommem[25382] <= 16'hD081;
rommem[25383] <= 16'h6900;
rommem[25384] <= 16'h023A;
rommem[25385] <= 16'h60EA;
rommem[25386] <= 16'h6100;
rommem[25387] <= 16'h044E;
rommem[25388] <= 16'h2D75;
rommem[25389] <= 16'h2F00;
rommem[25390] <= 16'h6100;
rommem[25391] <= 16'h000A;
rommem[25392] <= 16'h4480;
rommem[25393] <= 16'h4EF9;
rommem[25394] <= 16'hFFFC;
rommem[25395] <= 16'hC64A;
rommem[25396] <= 16'h6100;
rommem[25397] <= 16'h002C;
rommem[25398] <= 16'h6100;
rommem[25399] <= 16'h0436;
rommem[25400] <= 16'h2A0F;
rommem[25401] <= 16'h2F00;
rommem[25402] <= 16'h6100;
rommem[25403] <= 16'h0020;
rommem[25404] <= 16'h221F;
rommem[25405] <= 16'h6100;
rommem[25406] <= 16'h00A8;
rommem[25407] <= 16'h60EC;
rommem[25408] <= 16'h6100;
rommem[25409] <= 16'h0422;
rommem[25410] <= 16'h2F49;
rommem[25411] <= 16'h2F00;
rommem[25412] <= 16'h6100;
rommem[25413] <= 16'h000C;
rommem[25414] <= 16'h221F;
rommem[25415] <= 16'hC141;
rommem[25416] <= 16'h6100;
rommem[25417] <= 16'h00D4;
rommem[25418] <= 16'h60D6;
rommem[25419] <= 16'h43F9;
rommem[25420] <= 16'hFFFC;
rommem[25421] <= 16'hC14C;
rommem[25422] <= 16'h45F9;
rommem[25423] <= 16'hFFFC;
rommem[25424] <= 16'hC196;
rommem[25425] <= 16'h6000;
rommem[25426] <= 16'hFB1E;
rommem[25427] <= 16'h6100;
rommem[25428] <= 16'h002C;
rommem[25429] <= 16'h6508;
rommem[25430] <= 16'h2240;
rommem[25431] <= 16'h4280;
rommem[25432] <= 16'h2011;
rommem[25433] <= 16'h4E75;
rommem[25434] <= 16'h6100;
rommem[25435] <= 16'h0408;
rommem[25436] <= 16'h2001;
rommem[25437] <= 16'h4A82;
rommem[25438] <= 16'h66F4;
rommem[25439] <= 16'h6100;
rommem[25440] <= 16'h03E4;
rommem[25441] <= 16'h280D;
rommem[25442] <= 16'h6100;
rommem[25443] <= 16'hFEFC;
rommem[25444] <= 16'h6100;
rommem[25445] <= 16'h03DA;
rommem[25446] <= 16'h2903;
rommem[25447] <= 16'h4E75;
rommem[25448] <= 16'h6000;
rommem[25449] <= 16'h016C;
rommem[25450] <= 16'h6100;
rommem[25451] <= 16'h0420;
rommem[25452] <= 16'h4280;
rommem[25453] <= 16'h1010;
rommem[25454] <= 16'h0400;
rommem[25455] <= 16'h0040;
rommem[25456] <= 16'h6540;
rommem[25457] <= 16'h6628;
rommem[25458] <= 16'h5288;
rommem[25459] <= 16'h6100;
rommem[25460] <= 16'hFFD6;
rommem[25461] <= 16'hD080;
rommem[25462] <= 16'h6500;
rommem[25463] <= 16'h019C;
rommem[25464] <= 16'hD080;
rommem[25465] <= 16'h6500;
rommem[25466] <= 16'h0196;
rommem[25467] <= 16'h2F00;
rommem[25468] <= 16'h6100;
rommem[25469] <= 16'h00FA;
rommem[25470] <= 16'h221F;
rommem[25471] <= 16'hB081;
rommem[25472] <= 16'h6300;
rommem[25473] <= 16'h017E;
rommem[25474] <= 16'h2038;
rommem[25475] <= 16'h0628;
rommem[25476] <= 16'h9081;
rommem[25477] <= 16'h4E75;
rommem[25478] <= 16'hB03C;
rommem[25479] <= 16'h001B;
rommem[25480] <= 16'h0A3C;
rommem[25481] <= 16'h0001;
rommem[25482] <= 16'h650C;
rommem[25483] <= 16'h5288;
rommem[25484] <= 16'hD080;
rommem[25485] <= 16'hD080;
rommem[25486] <= 16'h2238;
rommem[25487] <= 16'h0628;
rommem[25488] <= 16'hD081;
rommem[25489] <= 16'h4E75;
rommem[25490] <= 16'h2801;
rommem[25491] <= 16'hB184;
rommem[25492] <= 16'h4A80;
rommem[25493] <= 16'h6A02;
rommem[25494] <= 16'h4480;
rommem[25495] <= 16'h4A81;
rommem[25496] <= 16'h6A02;
rommem[25497] <= 16'h4481;
rommem[25498] <= 16'hB2BC;
rommem[25499] <= 16'h0000;
rommem[25500] <= 16'hFFFF;
rommem[25501] <= 16'h630C;
rommem[25502] <= 16'hC141;
rommem[25503] <= 16'hB2BC;
rommem[25504] <= 16'h0000;
rommem[25505] <= 16'hFFFF;
rommem[25506] <= 16'h6200;
rommem[25507] <= 16'h0144;
rommem[25508] <= 16'h2400;
rommem[25509] <= 16'hC4C1;
rommem[25510] <= 16'h4840;
rommem[25511] <= 16'hC0C1;
rommem[25512] <= 16'h4840;
rommem[25513] <= 16'h4A80;
rommem[25514] <= 16'h6600;
rommem[25515] <= 16'h0134;
rommem[25516] <= 16'hD082;
rommem[25517] <= 16'h6B00;
rommem[25518] <= 16'h012E;
rommem[25519] <= 16'h4A84;
rommem[25520] <= 16'h6A02;
rommem[25521] <= 16'h4480;
rommem[25522] <= 16'h4E75;
rommem[25523] <= 16'h4A81;
rommem[25524] <= 16'h6700;
rommem[25525] <= 16'h0120;
rommem[25526] <= 16'h2401;
rommem[25527] <= 16'h2801;
rommem[25528] <= 16'hB184;
rommem[25529] <= 16'h4A80;
rommem[25530] <= 16'h6A02;
rommem[25531] <= 16'h4480;
rommem[25532] <= 16'h4A81;
rommem[25533] <= 16'h6A02;
rommem[25534] <= 16'h4481;
rommem[25535] <= 16'h761F;
rommem[25536] <= 16'h2200;
rommem[25537] <= 16'h4280;
rommem[25538] <= 16'hD281;
rommem[25539] <= 16'hD180;
rommem[25540] <= 16'h6708;
rommem[25541] <= 16'hB082;
rommem[25542] <= 16'h6B04;
rommem[25543] <= 16'h5281;
rommem[25544] <= 16'h9082;
rommem[25545] <= 16'h51CB;
rommem[25546] <= 16'hFFF0;
rommem[25547] <= 16'hC141;
rommem[25548] <= 16'h4A84;
rommem[25549] <= 16'h6A04;
rommem[25550] <= 16'h4480;
rommem[25551] <= 16'h4481;
rommem[25552] <= 16'h4E75;
rommem[25553] <= 16'h6100;
rommem[25554] <= 16'hFF1A;
rommem[25555] <= 16'h2240;
rommem[25556] <= 16'h4280;
rommem[25557] <= 16'h1011;
rommem[25558] <= 16'h4E75;
rommem[25559] <= 16'h6100;
rommem[25560] <= 16'hFF0E;
rommem[25561] <= 16'h4A80;
rommem[25562] <= 16'h6700;
rommem[25563] <= 16'h00D4;
rommem[25564] <= 16'h6B00;
rommem[25565] <= 16'h00D0;
rommem[25566] <= 16'h2200;
rommem[25567] <= 16'h2278;
rommem[25568] <= 16'h0600;
rommem[25569] <= 16'hB3FC;
rommem[25570] <= 16'hFFFC;
rommem[25571] <= 16'hCC5D;
rommem[25572] <= 16'h6506;
rommem[25573] <= 16'h43F9;
rommem[25574] <= 16'hFFFC;
rommem[25575] <= 16'hC000;
rommem[25576] <= 16'h2019;
rommem[25577] <= 16'h0880;
rommem[25578] <= 16'h001F;
rommem[25579] <= 16'h21C9;
rommem[25580] <= 16'h0600;
rommem[25581] <= 16'h6100;
rommem[25582] <= 16'hFF8A;
rommem[25583] <= 16'h2001;
rommem[25584] <= 16'h5280;
rommem[25585] <= 16'h4E75;
rommem[25586] <= 16'h6100;
rommem[25587] <= 16'hFED8;
rommem[25588] <= 16'h4A80;
rommem[25589] <= 16'h6A06;
rommem[25590] <= 16'h4480;
rommem[25591] <= 16'h6B00;
rommem[25592] <= 16'h009A;
rommem[25593] <= 16'h4E75;
rommem[25594] <= 16'h2038;
rommem[25595] <= 16'h0628;
rommem[25596] <= 16'h90B8;
rommem[25597] <= 16'h0624;
rommem[25598] <= 16'h4E75;
rommem[25599] <= 16'h6100;
rommem[25600] <= 16'hFED4;
rommem[25601] <= 16'h653A;
rommem[25602] <= 16'h2F00;
rommem[25603] <= 16'h6100;
rommem[25604] <= 16'h029C;
rommem[25605] <= 16'h3D0B;
rommem[25606] <= 16'h6100;
rommem[25607] <= 16'hFDB4;
rommem[25608] <= 16'h2C5F;
rommem[25609] <= 16'h2C80;
rommem[25610] <= 16'h4E75;
rommem[25611] <= 16'h6026;
rommem[25612] <= 16'h6100;
rommem[25613] <= 16'h028A;
rommem[25614] <= 16'h3A07;
rommem[25615] <= 16'h588F;
rommem[25616] <= 16'h6000;
rommem[25617] <= 16'hFA1C;
rommem[25618] <= 16'h6100;
rommem[25619] <= 16'h027E;
rommem[25620] <= 16'h0D07;
rommem[25621] <= 16'h588F;
rommem[25622] <= 16'h6000;
rommem[25623] <= 16'hF9F4;
rommem[25624] <= 16'h4E75;
rommem[25625] <= 16'h6100;
rommem[25626] <= 16'h02C2;
rommem[25627] <= 16'h0C10;
rommem[25628] <= 16'h000D;
rommem[25629] <= 16'h6602;
rommem[25630] <= 16'h4E75;
rommem[25631] <= 16'h2F08;
rommem[25632] <= 16'h4DF9;
rommem[25633] <= 16'hFFFC;
rommem[25634] <= 16'hCBDF;
rommem[25635] <= 16'h6100;
rommem[25636] <= 16'h031E;
rommem[25637] <= 16'h205F;
rommem[25638] <= 16'h2038;
rommem[25639] <= 16'h0604;
rommem[25640] <= 16'h6700;
rommem[25641] <= 16'hF80E;
rommem[25642] <= 16'hB0BC;
rommem[25643] <= 16'hFFFF;
rommem[25644] <= 16'hFFFF;
rommem[25645] <= 16'h6700;
rommem[25646] <= 16'hFBC2;
rommem[25647] <= 16'h1F10;
rommem[25648] <= 16'h4210;
rommem[25649] <= 16'h2278;
rommem[25650] <= 16'h0604;
rommem[25651] <= 16'h6100;
rommem[25652] <= 16'h0220;
rommem[25653] <= 16'h109F;
rommem[25654] <= 16'h103C;
rommem[25655] <= 16'h003F;
rommem[25656] <= 16'h6100;
rommem[25657] <= 16'hF796;
rommem[25658] <= 16'h4280;
rommem[25659] <= 16'h5389;
rommem[25660] <= 16'h6100;
rommem[25661] <= 16'h013E;
rommem[25662] <= 16'h6000;
rommem[25663] <= 16'hF7E2;
rommem[25664] <= 16'h2F08;
rommem[25665] <= 16'h4DF9;
rommem[25666] <= 16'hFFFC;
rommem[25667] <= 16'hCBE7;
rommem[25668] <= 16'h60BC;
rommem[25669] <= 16'h2F08;
rommem[25670] <= 16'h4DF9;
rommem[25671] <= 16'hFFFC;
rommem[25672] <= 16'hCBD8;
rommem[25673] <= 16'h60B2;
rommem[25674] <= 16'h6100;
rommem[25675] <= 16'hF772;
rommem[25676] <= 16'h103C;
rommem[25677] <= 16'h0020;
rommem[25678] <= 16'h6100;
rommem[25679] <= 16'hF76A;
rommem[25680] <= 16'h41F8;
rommem[25681] <= 16'h0630;
rommem[25682] <= 16'h6100;
rommem[25683] <= 16'h02A8;
rommem[25684] <= 16'h67FA;
rommem[25685] <= 16'hB03C;
rommem[25686] <= 16'h0008;
rommem[25687] <= 16'h6726;
rommem[25688] <= 16'hB03C;
rommem[25689] <= 16'h0018;
rommem[25690] <= 16'h6744;
rommem[25691] <= 16'hB03C;
rommem[25692] <= 16'h000D;
rommem[25693] <= 16'h6706;
rommem[25694] <= 16'hB03C;
rommem[25695] <= 16'h0020;
rommem[25696] <= 16'h65E2;
rommem[25697] <= 16'h10C0;
rommem[25698] <= 16'h6100;
rommem[25699] <= 16'hF742;
rommem[25700] <= 16'hB03C;
rommem[25701] <= 16'h000D;
rommem[25702] <= 16'h675C;
rommem[25703] <= 16'hB1FC;
rommem[25704] <= 16'h0000;
rommem[25705] <= 16'h067F;
rommem[25706] <= 16'h65CE;
rommem[25707] <= 16'h103C;
rommem[25708] <= 16'h0008;
rommem[25709] <= 16'h6100;
rommem[25710] <= 16'hF72C;
rommem[25711] <= 16'h103C;
rommem[25712] <= 16'h0020;
rommem[25713] <= 16'h6100;
rommem[25714] <= 16'hF724;
rommem[25715] <= 16'hB1FC;
rommem[25716] <= 16'h0000;
rommem[25717] <= 16'h0630;
rommem[25718] <= 16'h63B6;
rommem[25719] <= 16'h103C;
rommem[25720] <= 16'h0008;
rommem[25721] <= 16'h6100;
rommem[25722] <= 16'hF714;
rommem[25723] <= 16'h5388;
rommem[25724] <= 16'h60AA;
rommem[25725] <= 16'h2208;
rommem[25726] <= 16'h0481;
rommem[25727] <= 16'h0000;
rommem[25728] <= 16'h0630;
rommem[25729] <= 16'h671E;
rommem[25730] <= 16'h5381;
rommem[25731] <= 16'h103C;
rommem[25732] <= 16'h0008;
rommem[25733] <= 16'h6100;
rommem[25734] <= 16'hF6FC;
rommem[25735] <= 16'h103C;
rommem[25736] <= 16'h0020;
rommem[25737] <= 16'h6100;
rommem[25738] <= 16'hF6F4;
rommem[25739] <= 16'h103C;
rommem[25740] <= 16'h0008;
rommem[25741] <= 16'h6100;
rommem[25742] <= 16'hF6EC;
rommem[25743] <= 16'h51C9;
rommem[25744] <= 16'hFFE6;
rommem[25745] <= 16'h41F8;
rommem[25746] <= 16'h0630;
rommem[25747] <= 16'h6000;
rommem[25748] <= 16'hFF7C;
rommem[25749] <= 16'h103C;
rommem[25750] <= 16'h000A;
rommem[25751] <= 16'h6100;
rommem[25752] <= 16'hF6D8;
rommem[25753] <= 16'h4E75;
rommem[25754] <= 16'hB2BC;
rommem[25755] <= 16'h0000;
rommem[25756] <= 16'hFFFF;
rommem[25757] <= 16'h6400;
rommem[25758] <= 16'hFF4E;
rommem[25759] <= 16'h2279;
rommem[25760] <= 16'hFFFC;
rommem[25761] <= 16'hC01C;
rommem[25762] <= 16'h2478;
rommem[25763] <= 16'h0624;
rommem[25764] <= 16'h538A;
rommem[25765] <= 16'hB5C9;
rommem[25766] <= 16'h650C;
rommem[25767] <= 16'h1419;
rommem[25768] <= 16'hE18A;
rommem[25769] <= 16'h1411;
rommem[25770] <= 16'h5389;
rommem[25771] <= 16'hB481;
rommem[25772] <= 16'h6502;
rommem[25773] <= 16'h4E75;
rommem[25774] <= 16'h5489;
rommem[25775] <= 16'h0C19;
rommem[25776] <= 16'h000D;
rommem[25777] <= 16'h66FA;
rommem[25778] <= 16'h60DE;
rommem[25779] <= 16'hB7C9;
rommem[25780] <= 16'h6704;
rommem[25781] <= 16'h14D9;
rommem[25782] <= 16'h60F8;
rommem[25783] <= 16'h4E75;
rommem[25784] <= 16'hB5C9;
rommem[25785] <= 16'h67FA;
rommem[25786] <= 16'h1721;
rommem[25787] <= 16'h60F8;
rommem[25788] <= 16'h2C5F;
rommem[25789] <= 16'h21DF;
rommem[25790] <= 16'h0610;
rommem[25791] <= 16'h6710;
rommem[25792] <= 16'h21DF;
rommem[25793] <= 16'h0614;
rommem[25794] <= 16'h21DF;
rommem[25795] <= 16'h0618;
rommem[25796] <= 16'h21DF;
rommem[25797] <= 16'h061C;
rommem[25798] <= 16'h21DF;
rommem[25799] <= 16'h0620;
rommem[25800] <= 16'h4ED6;
rommem[25801] <= 16'h2238;
rommem[25802] <= 16'h062C;
rommem[25803] <= 16'h928F;
rommem[25804] <= 16'h6400;
rommem[25805] <= 16'hFEE6;
rommem[25806] <= 16'h2C5F;
rommem[25807] <= 16'h2238;
rommem[25808] <= 16'h0610;
rommem[25809] <= 16'h6710;
rommem[25810] <= 16'h2F38;
rommem[25811] <= 16'h0620;
rommem[25812] <= 16'h2F38;
rommem[25813] <= 16'h061C;
rommem[25814] <= 16'h2F38;
rommem[25815] <= 16'h0618;
rommem[25816] <= 16'h2F38;
rommem[25817] <= 16'h0614;
rommem[25818] <= 16'h2F01;
rommem[25819] <= 16'h4ED6;
rommem[25820] <= 16'h1200;
rommem[25821] <= 16'h1019;
rommem[25822] <= 16'hB200;
rommem[25823] <= 16'h6712;
rommem[25824] <= 16'h6100;
rommem[25825] <= 16'hF646;
rommem[25826] <= 16'hB03C;
rommem[25827] <= 16'h000D;
rommem[25828] <= 16'h66F0;
rommem[25829] <= 16'h103C;
rommem[25830] <= 16'h000A;
rommem[25831] <= 16'h6100;
rommem[25832] <= 16'hF638;
rommem[25833] <= 16'h4E75;
rommem[25834] <= 16'h6100;
rommem[25835] <= 16'h00CE;
rommem[25836] <= 16'h221B;
rommem[25837] <= 16'h103C;
rommem[25838] <= 16'h0022;
rommem[25839] <= 16'h2248;
rommem[25840] <= 16'h6100;
rommem[25841] <= 16'hFFD6;
rommem[25842] <= 16'h2049;
rommem[25843] <= 16'h225F;
rommem[25844] <= 16'hB03C;
rommem[25845] <= 16'h000A;
rommem[25846] <= 16'h6700;
rommem[25847] <= 16'hF834;
rommem[25848] <= 16'h5489;
rommem[25849] <= 16'h4ED1;
rommem[25850] <= 16'h6100;
rommem[25851] <= 16'h00AE;
rommem[25852] <= 16'h2707;
rommem[25853] <= 16'h103C;
rommem[25854] <= 16'h0027;
rommem[25855] <= 16'h60DE;
rommem[25856] <= 16'h6100;
rommem[25857] <= 16'h00A2;
rommem[25858] <= 16'h5F0D;
rommem[25859] <= 16'h103C;
rommem[25860] <= 16'h000D;
rommem[25861] <= 16'h6100;
rommem[25862] <= 16'hF5FC;
rommem[25863] <= 16'h225F;
rommem[25864] <= 16'h60DE;
rommem[25865] <= 16'h4E75;
rommem[25866] <= 16'h2601;
rommem[25867] <= 16'h2F04;
rommem[25868] <= 16'h1F3C;
rommem[25869] <= 16'h00FF;
rommem[25870] <= 16'h4A81;
rommem[25871] <= 16'h6A04;
rommem[25872] <= 16'h4481;
rommem[25873] <= 16'h5384;
rommem[25874] <= 16'h82FC;
rommem[25875] <= 16'h000A;
rommem[25876] <= 16'h690A;
rommem[25877] <= 16'h2001;
rommem[25878] <= 16'h0281;
rommem[25879] <= 16'h0000;
rommem[25880] <= 16'hFFFF;
rommem[25881] <= 16'h601A;
rommem[25882] <= 16'h2001;
rommem[25883] <= 16'h4241;
rommem[25884] <= 16'h4841;
rommem[25885] <= 16'h82FC;
rommem[25886] <= 16'h000A;
rommem[25887] <= 16'h2401;
rommem[25888] <= 16'h2200;
rommem[25889] <= 16'h82FC;
rommem[25890] <= 16'h000A;
rommem[25891] <= 16'h2001;
rommem[25892] <= 16'h4841;
rommem[25893] <= 16'h2202;
rommem[25894] <= 16'h4841;
rommem[25895] <= 16'h4840;
rommem[25896] <= 16'h1F00;
rommem[25897] <= 16'h4840;
rommem[25898] <= 16'h5384;
rommem[25899] <= 16'h4A81;
rommem[25900] <= 16'h66CA;
rommem[25901] <= 16'h5384;
rommem[25902] <= 16'h6B0C;
rommem[25903] <= 16'h103C;
rommem[25904] <= 16'h0020;
rommem[25905] <= 16'h6100;
rommem[25906] <= 16'hF5A4;
rommem[25907] <= 16'h51CC;
rommem[25908] <= 16'hFFF6;
rommem[25909] <= 16'h4A83;
rommem[25910] <= 16'h6A08;
rommem[25911] <= 16'h103C;
rommem[25912] <= 16'h002D;
rommem[25913] <= 16'h6100;
rommem[25914] <= 16'hF594;
rommem[25915] <= 16'h101F;
rommem[25916] <= 16'h6B0A;
rommem[25917] <= 16'h0600;
rommem[25918] <= 16'h0030;
rommem[25919] <= 16'h6100;
rommem[25920] <= 16'hF588;
rommem[25921] <= 16'h60F2;
rommem[25922] <= 16'h281F;
rommem[25923] <= 16'h4E75;
rommem[25924] <= 16'h4281;
rommem[25925] <= 16'h1219;
rommem[25926] <= 16'hE189;
rommem[25927] <= 16'h1219;
rommem[25928] <= 16'h7805;
rommem[25929] <= 16'h6100;
rommem[25930] <= 16'hFF80;
rommem[25931] <= 16'h103C;
rommem[25932] <= 16'h0020;
rommem[25933] <= 16'h6100;
rommem[25934] <= 16'hF56C;
rommem[25935] <= 16'h4280;
rommem[25936] <= 16'h6000;
rommem[25937] <= 16'hFF16;
rommem[25938] <= 16'h6100;
rommem[25939] <= 16'h0050;
rommem[25940] <= 16'h225F;
rommem[25941] <= 16'h1219;
rommem[25942] <= 16'hB210;
rommem[25943] <= 16'h6708;
rommem[25944] <= 16'h4281;
rommem[25945] <= 16'h1211;
rommem[25946] <= 16'hD3C1;
rommem[25947] <= 16'h4ED1;
rommem[25948] <= 16'h5288;
rommem[25949] <= 16'h5289;
rommem[25950] <= 16'h4ED1;
rommem[25951] <= 16'h4281;
rommem[25952] <= 16'h4282;
rommem[25953] <= 16'h6100;
rommem[25954] <= 16'h0032;
rommem[25955] <= 16'h0C10;
rommem[25956] <= 16'h0030;
rommem[25957] <= 16'h6528;
rommem[25958] <= 16'h0C10;
rommem[25959] <= 16'h0039;
rommem[25960] <= 16'h6222;
rommem[25961] <= 16'hB2BC;
rommem[25962] <= 16'h0CCC;
rommem[25963] <= 16'hCCCC;
rommem[25964] <= 16'h6400;
rommem[25965] <= 16'hFDB0;
rommem[25966] <= 16'h2001;
rommem[25967] <= 16'hD281;
rommem[25968] <= 16'hD281;
rommem[25969] <= 16'hD280;
rommem[25970] <= 16'hD281;
rommem[25971] <= 16'h1018;
rommem[25972] <= 16'h0280;
rommem[25973] <= 16'h0000;
rommem[25974] <= 16'h000F;
rommem[25975] <= 16'hD280;
rommem[25976] <= 16'h5282;
rommem[25977] <= 16'h60D2;
rommem[25978] <= 16'h4E75;
rommem[25979] <= 16'h0C10;
rommem[25980] <= 16'h0020;
rommem[25981] <= 16'h6604;
rommem[25982] <= 16'h5288;
rommem[25983] <= 16'h60F6;
rommem[25984] <= 16'h4E75;
rommem[25985] <= 16'h41F8;
rommem[25986] <= 16'h0630;
rommem[25987] <= 16'h4201;
rommem[25988] <= 16'h1018;
rommem[25989] <= 16'hB03C;
rommem[25990] <= 16'h000D;
rommem[25991] <= 16'h671A;
rommem[25992] <= 16'hB03C;
rommem[25993] <= 16'h0022;
rommem[25994] <= 16'h6716;
rommem[25995] <= 16'hB03C;
rommem[25996] <= 16'h0027;
rommem[25997] <= 16'h6710;
rommem[25998] <= 16'h4A01;
rommem[25999] <= 16'h66E8;
rommem[26000] <= 16'h6100;
rommem[26001] <= 16'h001A;
rommem[26002] <= 16'h1100;
rommem[26003] <= 16'h5288;
rommem[26004] <= 16'h60DE;
rommem[26005] <= 16'h4E75;
rommem[26006] <= 16'h4A01;
rommem[26007] <= 16'h6604;
rommem[26008] <= 16'h1200;
rommem[26009] <= 16'h60D4;
rommem[26010] <= 16'hB200;
rommem[26011] <= 16'h66D0;
rommem[26012] <= 16'h4201;
rommem[26013] <= 16'h60CC;
rommem[26014] <= 16'hB03C;
rommem[26015] <= 16'h0061;
rommem[26016] <= 16'h650A;
rommem[26017] <= 16'hB03C;
rommem[26018] <= 16'h007A;
rommem[26019] <= 16'h6204;
rommem[26020] <= 16'h0400;
rommem[26021] <= 16'h0020;
rommem[26022] <= 16'h4E75;
rommem[26023] <= 16'h6100;
rommem[26024] <= 16'hF4BC;
rommem[26025] <= 16'h670A;
rommem[26026] <= 16'hB03C;
rommem[26027] <= 16'h0003;
rommem[26028] <= 16'h6604;
rommem[26029] <= 16'h6000;
rommem[26030] <= 16'hF504;
rommem[26031] <= 16'h4E75;
rommem[26032] <= 16'h4DF9;
rommem[26033] <= 16'hFFFC;
rommem[26034] <= 16'hCBED;
rommem[26035] <= 16'h101E;
rommem[26036] <= 16'h6706;
rommem[26037] <= 16'h6100;
rommem[26038] <= 16'hF49C;
rommem[26039] <= 16'h60F6;
rommem[26040] <= 16'h4E75;
rommem[26041] <= 16'h48E7;
rommem[26042] <= 16'hC000;
rommem[26043] <= 16'h2200;
rommem[26044] <= 16'h7006;
rommem[26045] <= 16'h4E4F;
rommem[26046] <= 16'h4CDF;
rommem[26047] <= 16'h0003;
rommem[26048] <= 16'h4E75;
rommem[26049] <= 16'h2F01;
rommem[26050] <= 16'h7007;
rommem[26051] <= 16'h4E4F;
rommem[26052] <= 16'h4A00;
rommem[26053] <= 16'h670A;
rommem[26054] <= 16'h7005;
rommem[26055] <= 16'h4E4F;
rommem[26056] <= 16'h2001;
rommem[26057] <= 16'h221F;
rommem[26058] <= 16'h4A00;
rommem[26059] <= 16'h4E75;
rommem[26060] <= 16'h0839;
rommem[26061] <= 16'h0005;
rommem[26062] <= 16'hFFDC;
rommem[26063] <= 16'h0A01;
rommem[26064] <= 16'h67F6;
rommem[26065] <= 16'h13C0;
rommem[26066] <= 16'hFFDC;
rommem[26067] <= 16'h0A00;
rommem[26068] <= 16'h4E75;
rommem[26069] <= 16'h0839;
rommem[26070] <= 16'h0000;
rommem[26071] <= 16'hFFDC;
rommem[26072] <= 16'h0A01;
rommem[26073] <= 16'h670A;
rommem[26074] <= 16'h1039;
rommem[26075] <= 16'hFFDC;
rommem[26076] <= 16'h0A00;
rommem[26077] <= 16'h0200;
rommem[26078] <= 16'h007F;
rommem[26079] <= 16'h4E75;
rommem[26080] <= 16'h1E3C;
rommem[26081] <= 16'h00E4;
rommem[26082] <= 16'h4E4E;
rommem[26083] <= 16'h0D0A;
rommem[26084] <= 16'h476F;
rommem[26085] <= 16'h7264;
rommem[26086] <= 16'h6F0D;
rommem[26087] <= 16'h0A0A;
rommem[26088] <= 16'h000D;
rommem[26089] <= 16'h0A4F;
rommem[26090] <= 16'h4B0D;
rommem[26091] <= 16'h0A00;
rommem[26092] <= 16'h486F;
rommem[26093] <= 16'h773F;
rommem[26094] <= 16'h0D0A;
rommem[26095] <= 16'h0057;
rommem[26096] <= 16'h6861;
rommem[26097] <= 16'h743F;
rommem[26098] <= 16'h0D0A;
rommem[26099] <= 16'h0053;
rommem[26100] <= 16'h6F72;
rommem[26101] <= 16'h7279;
rommem[26102] <= 16'h2E0D;
rommem[26103] <= 16'h0A00;
