// ============================================================================
//        __
//   \\__/ o\    (C) 2020  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	div_lut.sv
//    - divide reciprocal lookup table
//    - 2048 entries (1 block ram)
//
//
// This source file is free software: you can redistribute it and/or modify 
// it under the terms of the GNU Lesser General Public License as published 
// by the Free Software Foundation, either version 3 of the License, or     
// (at your option) any later version.                                      
//                                                                          
// This source file is distributed in the hope that it will be useful,      
// but WITHOUT ANY WARRANTY; without even the implied warranty of           
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the            
// GNU General Public License for more details.                             
//                                                                          
// You should have received a copy of the GNU General Public License        
// along with this program.  If not, see <http://www.gnu.org/licenses/>.    
//                                                                          
// ============================================================================

module div_lut(clk, ce, i, o);
input clk;
input ce;
input [10:0] i;
output reg [15:0] o;

always @(posedge clk)
if (ce)
case(i)
11'h000: o <= 16'hFFFF;
11'h001: o <= 16'hFFE0;
11'h002: o <= 16'hFFC0;
11'h003: o <= 16'hFFA0;
11'h004: o <= 16'hFF80;
11'h005: o <= 16'hFF60;
11'h006: o <= 16'hFF40;
11'h007: o <= 16'hFF20;
11'h008: o <= 16'hFF00;
11'h009: o <= 16'hFEE1;
11'h00A: o <= 16'hFEC1;
11'h00B: o <= 16'hFEA1;
11'h00C: o <= 16'hFE82;
11'h00D: o <= 16'hFE62;
11'h00E: o <= 16'hFE43;
11'h00F: o <= 16'hFE23;
11'h010: o <= 16'hFE03;
11'h011: o <= 16'hFDE4;
11'h012: o <= 16'hFDC5;
11'h013: o <= 16'hFDA5;
11'h014: o <= 16'hFD86;
11'h015: o <= 16'hFD66;
11'h016: o <= 16'hFD47;
11'h017: o <= 16'hFD28;
11'h018: o <= 16'hFD08;
11'h019: o <= 16'hFCE9;
11'h01A: o <= 16'hFCCA;
11'h01B: o <= 16'hFCAB;
11'h01C: o <= 16'hFC8C;
11'h01D: o <= 16'hFC6C;
11'h01E: o <= 16'hFC4D;
11'h01F: o <= 16'hFC2E;
11'h020: o <= 16'hFC0F;
11'h021: o <= 16'hFBF0;
11'h022: o <= 16'hFBD1;
11'h023: o <= 16'hFBB2;
11'h024: o <= 16'hFB93;
11'h025: o <= 16'hFB75;
11'h026: o <= 16'hFB56;
11'h027: o <= 16'hFB37;
11'h028: o <= 16'hFB18;
11'h029: o <= 16'hFAF9;
11'h02A: o <= 16'hFADB;
11'h02B: o <= 16'hFABC;
11'h02C: o <= 16'hFA9D;
11'h02D: o <= 16'hFA7E;
11'h02E: o <= 16'hFA60;
11'h02F: o <= 16'hFA41;
11'h030: o <= 16'hFA23;
11'h031: o <= 16'hFA04;
11'h032: o <= 16'hF9E6;
11'h033: o <= 16'hF9C7;
11'h034: o <= 16'hF9A9;
11'h035: o <= 16'hF98A;
11'h036: o <= 16'hF96C;
11'h037: o <= 16'hF94E;
11'h038: o <= 16'hF92F;
11'h039: o <= 16'hF911;
11'h03A: o <= 16'hF8F3;
11'h03B: o <= 16'hF8D4;
11'h03C: o <= 16'hF8B6;
11'h03D: o <= 16'hF898;
11'h03E: o <= 16'hF87A;
11'h03F: o <= 16'hF85C;
11'h040: o <= 16'hF83E;
11'h041: o <= 16'hF81F;
11'h042: o <= 16'hF801;
11'h043: o <= 16'hF7E3;
11'h044: o <= 16'hF7C5;
11'h045: o <= 16'hF7A7;
11'h046: o <= 16'hF78A;
11'h047: o <= 16'hF76C;
11'h048: o <= 16'hF74E;
11'h049: o <= 16'hF730;
11'h04A: o <= 16'hF712;
11'h04B: o <= 16'hF6F4;
11'h04C: o <= 16'hF6D7;
11'h04D: o <= 16'hF6B9;
11'h04E: o <= 16'hF69B;
11'h04F: o <= 16'hF67D;
11'h050: o <= 16'hF660;
11'h051: o <= 16'hF642;
11'h052: o <= 16'hF625;
11'h053: o <= 16'hF607;
11'h054: o <= 16'hF5E9;
11'h055: o <= 16'hF5CC;
11'h056: o <= 16'hF5AE;
11'h057: o <= 16'hF591;
11'h058: o <= 16'hF574;
11'h059: o <= 16'hF556;
11'h05A: o <= 16'hF539;
11'h05B: o <= 16'hF51B;
11'h05C: o <= 16'hF4FE;
11'h05D: o <= 16'hF4E1;
11'h05E: o <= 16'hF4C4;
11'h05F: o <= 16'hF4A6;
11'h060: o <= 16'hF489;
11'h061: o <= 16'hF46C;
11'h062: o <= 16'hF44F;
11'h063: o <= 16'hF432;
11'h064: o <= 16'hF414;
11'h065: o <= 16'hF3F7;
11'h066: o <= 16'hF3DA;
11'h067: o <= 16'hF3BD;
11'h068: o <= 16'hF3A0;
11'h069: o <= 16'hF383;
11'h06A: o <= 16'hF366;
11'h06B: o <= 16'hF34A;
11'h06C: o <= 16'hF32D;
11'h06D: o <= 16'hF310;
11'h06E: o <= 16'hF2F3;
11'h06F: o <= 16'hF2D6;
11'h070: o <= 16'hF2B9;
11'h071: o <= 16'hF29D;
11'h072: o <= 16'hF280;
11'h073: o <= 16'hF263;
11'h074: o <= 16'hF246;
11'h075: o <= 16'hF22A;
11'h076: o <= 16'hF20D;
11'h077: o <= 16'hF1F1;
11'h078: o <= 16'hF1D4;
11'h079: o <= 16'hF1B8;
11'h07A: o <= 16'hF19B;
11'h07B: o <= 16'hF17E;
11'h07C: o <= 16'hF162;
11'h07D: o <= 16'hF146;
11'h07E: o <= 16'hF129;
11'h07F: o <= 16'hF10D;
11'h080: o <= 16'hF0F0;
11'h081: o <= 16'hF0D4;
11'h082: o <= 16'hF0B8;
11'h083: o <= 16'hF09C;
11'h084: o <= 16'hF07F;
11'h085: o <= 16'hF063;
11'h086: o <= 16'hF047;
11'h087: o <= 16'hF02B;
11'h088: o <= 16'hF00F;
11'h089: o <= 16'hEFF2;
11'h08A: o <= 16'hEFD6;
11'h08B: o <= 16'hEFBA;
11'h08C: o <= 16'hEF9E;
11'h08D: o <= 16'hEF82;
11'h08E: o <= 16'hEF66;
11'h08F: o <= 16'hEF4A;
11'h090: o <= 16'hEF2E;
11'h091: o <= 16'hEF12;
11'h092: o <= 16'hEEF6;
11'h093: o <= 16'hEEDB;
11'h094: o <= 16'hEEBF;
11'h095: o <= 16'hEEA3;
11'h096: o <= 16'hEE87;
11'h097: o <= 16'hEE6B;
11'h098: o <= 16'hEE50;
11'h099: o <= 16'hEE34;
11'h09A: o <= 16'hEE18;
11'h09B: o <= 16'hEDFC;
11'h09C: o <= 16'hEDE1;
11'h09D: o <= 16'hEDC5;
11'h09E: o <= 16'hEDAA;
11'h09F: o <= 16'hED8E;
11'h0A0: o <= 16'hED73;
11'h0A1: o <= 16'hED57;
11'h0A2: o <= 16'hED3C;
11'h0A3: o <= 16'hED20;
11'h0A4: o <= 16'hED05;
11'h0A5: o <= 16'hECE9;
11'h0A6: o <= 16'hECCE;
11'h0A7: o <= 16'hECB2;
11'h0A8: o <= 16'hEC97;
11'h0A9: o <= 16'hEC7C;
11'h0AA: o <= 16'hEC60;
11'h0AB: o <= 16'hEC45;
11'h0AC: o <= 16'hEC2A;
11'h0AD: o <= 16'hEC0F;
11'h0AE: o <= 16'hEBF4;
11'h0AF: o <= 16'hEBD8;
11'h0B0: o <= 16'hEBBD;
11'h0B1: o <= 16'hEBA2;
11'h0B2: o <= 16'hEB87;
11'h0B3: o <= 16'hEB6C;
11'h0B4: o <= 16'hEB51;
11'h0B5: o <= 16'hEB36;
11'h0B6: o <= 16'hEB1B;
11'h0B7: o <= 16'hEB00;
11'h0B8: o <= 16'hEAE5;
11'h0B9: o <= 16'hEACA;
11'h0BA: o <= 16'hEAAF;
11'h0BB: o <= 16'hEA94;
11'h0BC: o <= 16'hEA79;
11'h0BD: o <= 16'hEA5E;
11'h0BE: o <= 16'hEA44;
11'h0BF: o <= 16'hEA29;
11'h0C0: o <= 16'hEA0E;
11'h0C1: o <= 16'hE9F3;
11'h0C2: o <= 16'hE9D9;
11'h0C3: o <= 16'hE9BE;
11'h0C4: o <= 16'hE9A3;
11'h0C5: o <= 16'hE989;
11'h0C6: o <= 16'hE96E;
11'h0C7: o <= 16'hE953;
11'h0C8: o <= 16'hE939;
11'h0C9: o <= 16'hE91E;
11'h0CA: o <= 16'hE904;
11'h0CB: o <= 16'hE8E9;
11'h0CC: o <= 16'hE8CF;
11'h0CD: o <= 16'hE8B4;
11'h0CE: o <= 16'hE89A;
11'h0CF: o <= 16'hE880;
11'h0D0: o <= 16'hE865;
11'h0D1: o <= 16'hE84B;
11'h0D2: o <= 16'hE830;
11'h0D3: o <= 16'hE816;
11'h0D4: o <= 16'hE7FC;
11'h0D5: o <= 16'hE7E2;
11'h0D6: o <= 16'hE7C7;
11'h0D7: o <= 16'hE7AD;
11'h0D8: o <= 16'hE793;
11'h0D9: o <= 16'hE779;
11'h0DA: o <= 16'hE75F;
11'h0DB: o <= 16'hE744;
11'h0DC: o <= 16'hE72A;
11'h0DD: o <= 16'hE710;
11'h0DE: o <= 16'hE6F6;
11'h0DF: o <= 16'hE6DC;
11'h0E0: o <= 16'hE6C2;
11'h0E1: o <= 16'hE6A8;
11'h0E2: o <= 16'hE68E;
11'h0E3: o <= 16'hE674;
11'h0E4: o <= 16'hE65A;
11'h0E5: o <= 16'hE640;
11'h0E6: o <= 16'hE627;
11'h0E7: o <= 16'hE60D;
11'h0E8: o <= 16'hE5F3;
11'h0E9: o <= 16'hE5D9;
11'h0EA: o <= 16'hE5BF;
11'h0EB: o <= 16'hE5A6;
11'h0EC: o <= 16'hE58C;
11'h0ED: o <= 16'hE572;
11'h0EE: o <= 16'hE558;
11'h0EF: o <= 16'hE53F;
11'h0F0: o <= 16'hE525;
11'h0F1: o <= 16'hE50B;
11'h0F2: o <= 16'hE4F2;
11'h0F3: o <= 16'hE4D8;
11'h0F4: o <= 16'hE4BF;
11'h0F5: o <= 16'hE4A5;
11'h0F6: o <= 16'hE48C;
11'h0F7: o <= 16'hE472;
11'h0F8: o <= 16'hE459;
11'h0F9: o <= 16'hE43F;
11'h0FA: o <= 16'hE426;
11'h0FB: o <= 16'hE40C;
11'h0FC: o <= 16'hE3F3;
11'h0FD: o <= 16'hE3DA;
11'h0FE: o <= 16'hE3C0;
11'h0FF: o <= 16'hE3A7;
11'h100: o <= 16'hE38E;
11'h101: o <= 16'hE374;
11'h102: o <= 16'hE35B;
11'h103: o <= 16'hE342;
11'h104: o <= 16'hE329;
11'h105: o <= 16'hE310;
11'h106: o <= 16'hE2F6;
11'h107: o <= 16'hE2DD;
11'h108: o <= 16'hE2C4;
11'h109: o <= 16'hE2AB;
11'h10A: o <= 16'hE292;
11'h10B: o <= 16'hE279;
11'h10C: o <= 16'hE260;
11'h10D: o <= 16'hE247;
11'h10E: o <= 16'hE22E;
11'h10F: o <= 16'hE215;
11'h110: o <= 16'hE1FC;
11'h111: o <= 16'hE1E3;
11'h112: o <= 16'hE1CA;
11'h113: o <= 16'hE1B1;
11'h114: o <= 16'hE198;
11'h115: o <= 16'hE180;
11'h116: o <= 16'hE167;
11'h117: o <= 16'hE14E;
11'h118: o <= 16'hE135;
11'h119: o <= 16'hE11C;
11'h11A: o <= 16'hE104;
11'h11B: o <= 16'hE0EB;
11'h11C: o <= 16'hE0D2;
11'h11D: o <= 16'hE0BA;
11'h11E: o <= 16'hE0A1;
11'h11F: o <= 16'hE088;
11'h120: o <= 16'hE070;
11'h121: o <= 16'hE057;
11'h122: o <= 16'hE03F;
11'h123: o <= 16'hE026;
11'h124: o <= 16'hE00E;
11'h125: o <= 16'hDFF5;
11'h126: o <= 16'hDFDD;
11'h127: o <= 16'hDFC4;
11'h128: o <= 16'hDFAC;
11'h129: o <= 16'hDF93;
11'h12A: o <= 16'hDF7B;
11'h12B: o <= 16'hDF62;
11'h12C: o <= 16'hDF4A;
11'h12D: o <= 16'hDF32;
11'h12E: o <= 16'hDF19;
11'h12F: o <= 16'hDF01;
11'h130: o <= 16'hDEE9;
11'h131: o <= 16'hDED1;
11'h132: o <= 16'hDEB8;
11'h133: o <= 16'hDEA0;
11'h134: o <= 16'hDE88;
11'h135: o <= 16'hDE70;
11'h136: o <= 16'hDE58;
11'h137: o <= 16'hDE40;
11'h138: o <= 16'hDE27;
11'h139: o <= 16'hDE0F;
11'h13A: o <= 16'hDDF7;
11'h13B: o <= 16'hDDDF;
11'h13C: o <= 16'hDDC7;
11'h13D: o <= 16'hDDAF;
11'h13E: o <= 16'hDD97;
11'h13F: o <= 16'hDD7F;
11'h140: o <= 16'hDD67;
11'h141: o <= 16'hDD4F;
11'h142: o <= 16'hDD37;
11'h143: o <= 16'hDD20;
11'h144: o <= 16'hDD08;
11'h145: o <= 16'hDCF0;
11'h146: o <= 16'hDCD8;
11'h147: o <= 16'hDCC0;
11'h148: o <= 16'hDCA8;
11'h149: o <= 16'hDC91;
11'h14A: o <= 16'hDC79;
11'h14B: o <= 16'hDC61;
11'h14C: o <= 16'hDC4A;
11'h14D: o <= 16'hDC32;
11'h14E: o <= 16'hDC1A;
11'h14F: o <= 16'hDC03;
11'h150: o <= 16'hDBEB;
11'h151: o <= 16'hDBD3;
11'h152: o <= 16'hDBBC;
11'h153: o <= 16'hDBA4;
11'h154: o <= 16'hDB8D;
11'h155: o <= 16'hDB75;
11'h156: o <= 16'hDB5E;
11'h157: o <= 16'hDB46;
11'h158: o <= 16'hDB2F;
11'h159: o <= 16'hDB17;
11'h15A: o <= 16'hDB00;
11'h15B: o <= 16'hDAE8;
11'h15C: o <= 16'hDAD1;
11'h15D: o <= 16'hDABA;
11'h15E: o <= 16'hDAA2;
11'h15F: o <= 16'hDA8B;
11'h160: o <= 16'hDA74;
11'h161: o <= 16'hDA5C;
11'h162: o <= 16'hDA45;
11'h163: o <= 16'hDA2E;
11'h164: o <= 16'hDA17;
11'h165: o <= 16'hD9FF;
11'h166: o <= 16'hD9E8;
11'h167: o <= 16'hD9D1;
11'h168: o <= 16'hD9BA;
11'h169: o <= 16'hD9A3;
11'h16A: o <= 16'hD98C;
11'h16B: o <= 16'hD974;
11'h16C: o <= 16'hD95D;
11'h16D: o <= 16'hD946;
11'h16E: o <= 16'hD92F;
11'h16F: o <= 16'hD918;
11'h170: o <= 16'hD901;
11'h171: o <= 16'hD8EA;
11'h172: o <= 16'hD8D3;
11'h173: o <= 16'hD8BC;
11'h174: o <= 16'hD8A5;
11'h175: o <= 16'hD88E;
11'h176: o <= 16'hD878;
11'h177: o <= 16'hD861;
11'h178: o <= 16'hD84A;
11'h179: o <= 16'hD833;
11'h17A: o <= 16'hD81C;
11'h17B: o <= 16'hD805;
11'h17C: o <= 16'hD7EF;
11'h17D: o <= 16'hD7D8;
11'h17E: o <= 16'hD7C1;
11'h17F: o <= 16'hD7AA;
11'h180: o <= 16'hD794;
11'h181: o <= 16'hD77D;
11'h182: o <= 16'hD766;
11'h183: o <= 16'hD750;
11'h184: o <= 16'hD739;
11'h185: o <= 16'hD722;
11'h186: o <= 16'hD70C;
11'h187: o <= 16'hD6F5;
11'h188: o <= 16'hD6DF;
11'h189: o <= 16'hD6C8;
11'h18A: o <= 16'hD6B2;
11'h18B: o <= 16'hD69B;
11'h18C: o <= 16'hD685;
11'h18D: o <= 16'hD66E;
11'h18E: o <= 16'hD658;
11'h18F: o <= 16'hD641;
11'h190: o <= 16'hD62B;
11'h191: o <= 16'hD615;
11'h192: o <= 16'hD5FE;
11'h193: o <= 16'hD5E8;
11'h194: o <= 16'hD5D2;
11'h195: o <= 16'hD5BB;
11'h196: o <= 16'hD5A5;
11'h197: o <= 16'hD58F;
11'h198: o <= 16'hD578;
11'h199: o <= 16'hD562;
11'h19A: o <= 16'hD54C;
11'h19B: o <= 16'hD536;
11'h19C: o <= 16'hD520;
11'h19D: o <= 16'hD509;
11'h19E: o <= 16'hD4F3;
11'h19F: o <= 16'hD4DD;
11'h1A0: o <= 16'hD4C7;
11'h1A1: o <= 16'hD4B1;
11'h1A2: o <= 16'hD49B;
11'h1A3: o <= 16'hD485;
11'h1A4: o <= 16'hD46F;
11'h1A5: o <= 16'hD459;
11'h1A6: o <= 16'hD443;
11'h1A7: o <= 16'hD42D;
11'h1A8: o <= 16'hD417;
11'h1A9: o <= 16'hD401;
11'h1AA: o <= 16'hD3EB;
11'h1AB: o <= 16'hD3D5;
11'h1AC: o <= 16'hD3BF;
11'h1AD: o <= 16'hD3A9;
11'h1AE: o <= 16'hD393;
11'h1AF: o <= 16'hD37D;
11'h1B0: o <= 16'hD368;
11'h1B1: o <= 16'hD352;
11'h1B2: o <= 16'hD33C;
11'h1B3: o <= 16'hD326;
11'h1B4: o <= 16'hD310;
11'h1B5: o <= 16'hD2FB;
11'h1B6: o <= 16'hD2E5;
11'h1B7: o <= 16'hD2CF;
11'h1B8: o <= 16'hD2BA;
11'h1B9: o <= 16'hD2A4;
11'h1BA: o <= 16'hD28E;
11'h1BB: o <= 16'hD279;
11'h1BC: o <= 16'hD263;
11'h1BD: o <= 16'hD24D;
11'h1BE: o <= 16'hD238;
11'h1BF: o <= 16'hD222;
11'h1C0: o <= 16'hD20D;
11'h1C1: o <= 16'hD1F7;
11'h1C2: o <= 16'hD1E2;
11'h1C3: o <= 16'hD1CC;
11'h1C4: o <= 16'hD1B7;
11'h1C5: o <= 16'hD1A1;
11'h1C6: o <= 16'hD18C;
11'h1C7: o <= 16'hD176;
11'h1C8: o <= 16'hD161;
11'h1C9: o <= 16'hD14B;
11'h1CA: o <= 16'hD136;
11'h1CB: o <= 16'hD121;
11'h1CC: o <= 16'hD10B;
11'h1CD: o <= 16'hD0F6;
11'h1CE: o <= 16'hD0E1;
11'h1CF: o <= 16'hD0CB;
11'h1D0: o <= 16'hD0B6;
11'h1D1: o <= 16'hD0A1;
11'h1D2: o <= 16'hD08C;
11'h1D3: o <= 16'hD076;
11'h1D4: o <= 16'hD061;
11'h1D5: o <= 16'hD04C;
11'h1D6: o <= 16'hD037;
11'h1D7: o <= 16'hD022;
11'h1D8: o <= 16'hD00D;
11'h1D9: o <= 16'hCFF7;
11'h1DA: o <= 16'hCFE2;
11'h1DB: o <= 16'hCFCD;
11'h1DC: o <= 16'hCFB8;
11'h1DD: o <= 16'hCFA3;
11'h1DE: o <= 16'hCF8E;
11'h1DF: o <= 16'hCF79;
11'h1E0: o <= 16'hCF64;
11'h1E1: o <= 16'hCF4F;
11'h1E2: o <= 16'hCF3A;
11'h1E3: o <= 16'hCF25;
11'h1E4: o <= 16'hCF10;
11'h1E5: o <= 16'hCEFB;
11'h1E6: o <= 16'hCEE6;
11'h1E7: o <= 16'hCED1;
11'h1E8: o <= 16'hCEBC;
11'h1E9: o <= 16'hCEA8;
11'h1EA: o <= 16'hCE93;
11'h1EB: o <= 16'hCE7E;
11'h1EC: o <= 16'hCE69;
11'h1ED: o <= 16'hCE54;
11'h1EE: o <= 16'hCE40;
11'h1EF: o <= 16'hCE2B;
11'h1F0: o <= 16'hCE16;
11'h1F1: o <= 16'hCE01;
11'h1F2: o <= 16'hCDED;
11'h1F3: o <= 16'hCDD8;
11'h1F4: o <= 16'hCDC3;
11'h1F5: o <= 16'hCDAF;
11'h1F6: o <= 16'hCD9A;
11'h1F7: o <= 16'hCD85;
11'h1F8: o <= 16'hCD71;
11'h1F9: o <= 16'hCD5C;
11'h1FA: o <= 16'hCD47;
11'h1FB: o <= 16'hCD33;
11'h1FC: o <= 16'hCD1E;
11'h1FD: o <= 16'hCD0A;
11'h1FE: o <= 16'hCCF5;
11'h1FF: o <= 16'hCCE1;
11'h200: o <= 16'hCCCC;
11'h201: o <= 16'hCCB8;
11'h202: o <= 16'hCCA3;
11'h203: o <= 16'hCC8F;
11'h204: o <= 16'hCC7B;
11'h205: o <= 16'hCC66;
11'h206: o <= 16'hCC52;
11'h207: o <= 16'hCC3D;
11'h208: o <= 16'hCC29;
11'h209: o <= 16'hCC15;
11'h20A: o <= 16'hCC00;
11'h20B: o <= 16'hCBEC;
11'h20C: o <= 16'hCBD8;
11'h20D: o <= 16'hCBC3;
11'h20E: o <= 16'hCBAF;
11'h20F: o <= 16'hCB9B;
11'h210: o <= 16'hCB87;
11'h211: o <= 16'hCB72;
11'h212: o <= 16'hCB5E;
11'h213: o <= 16'hCB4A;
11'h214: o <= 16'hCB36;
11'h215: o <= 16'hCB22;
11'h216: o <= 16'hCB0E;
11'h217: o <= 16'hCAF9;
11'h218: o <= 16'hCAE5;
11'h219: o <= 16'hCAD1;
11'h21A: o <= 16'hCABD;
11'h21B: o <= 16'hCAA9;
11'h21C: o <= 16'hCA95;
11'h21D: o <= 16'hCA81;
11'h21E: o <= 16'hCA6D;
11'h21F: o <= 16'hCA59;
11'h220: o <= 16'hCA45;
11'h221: o <= 16'hCA31;
11'h222: o <= 16'hCA1D;
11'h223: o <= 16'hCA09;
11'h224: o <= 16'hC9F5;
11'h225: o <= 16'hC9E1;
11'h226: o <= 16'hC9CD;
11'h227: o <= 16'hC9BA;
11'h228: o <= 16'hC9A6;
11'h229: o <= 16'hC992;
11'h22A: o <= 16'hC97E;
11'h22B: o <= 16'hC96A;
11'h22C: o <= 16'hC956;
11'h22D: o <= 16'hC943;
11'h22E: o <= 16'hC92F;
11'h22F: o <= 16'hC91B;
11'h230: o <= 16'hC907;
11'h231: o <= 16'hC8F4;
11'h232: o <= 16'hC8E0;
11'h233: o <= 16'hC8CC;
11'h234: o <= 16'hC8B9;
11'h235: o <= 16'hC8A5;
11'h236: o <= 16'hC891;
11'h237: o <= 16'hC87E;
11'h238: o <= 16'hC86A;
11'h239: o <= 16'hC856;
11'h23A: o <= 16'hC843;
11'h23B: o <= 16'hC82F;
11'h23C: o <= 16'hC81C;
11'h23D: o <= 16'hC808;
11'h23E: o <= 16'hC7F5;
11'h23F: o <= 16'hC7E1;
11'h240: o <= 16'hC7CE;
11'h241: o <= 16'hC7BA;
11'h242: o <= 16'hC7A7;
11'h243: o <= 16'hC793;
11'h244: o <= 16'hC780;
11'h245: o <= 16'hC76C;
11'h246: o <= 16'hC759;
11'h247: o <= 16'hC745;
11'h248: o <= 16'hC732;
11'h249: o <= 16'hC71F;
11'h24A: o <= 16'hC70B;
11'h24B: o <= 16'hC6F8;
11'h24C: o <= 16'hC6E5;
11'h24D: o <= 16'hC6D1;
11'h24E: o <= 16'hC6BE;
11'h24F: o <= 16'hC6AB;
11'h250: o <= 16'hC698;
11'h251: o <= 16'hC684;
11'h252: o <= 16'hC671;
11'h253: o <= 16'hC65E;
11'h254: o <= 16'hC64B;
11'h255: o <= 16'hC637;
11'h256: o <= 16'hC624;
11'h257: o <= 16'hC611;
11'h258: o <= 16'hC5FE;
11'h259: o <= 16'hC5EB;
11'h25A: o <= 16'hC5D8;
11'h25B: o <= 16'hC5C5;
11'h25C: o <= 16'hC5B2;
11'h25D: o <= 16'hC59E;
11'h25E: o <= 16'hC58B;
11'h25F: o <= 16'hC578;
11'h260: o <= 16'hC565;
11'h261: o <= 16'hC552;
11'h262: o <= 16'hC53F;
11'h263: o <= 16'hC52C;
11'h264: o <= 16'hC519;
11'h265: o <= 16'hC506;
11'h266: o <= 16'hC4F3;
11'h267: o <= 16'hC4E0;
11'h268: o <= 16'hC4CE;
11'h269: o <= 16'hC4BB;
11'h26A: o <= 16'hC4A8;
11'h26B: o <= 16'hC495;
11'h26C: o <= 16'hC482;
11'h26D: o <= 16'hC46F;
11'h26E: o <= 16'hC45C;
11'h26F: o <= 16'hC449;
11'h270: o <= 16'hC437;
11'h271: o <= 16'hC424;
11'h272: o <= 16'hC411;
11'h273: o <= 16'hC3FE;
11'h274: o <= 16'hC3EC;
11'h275: o <= 16'hC3D9;
11'h276: o <= 16'hC3C6;
11'h277: o <= 16'hC3B3;
11'h278: o <= 16'hC3A1;
11'h279: o <= 16'hC38E;
11'h27A: o <= 16'hC37B;
11'h27B: o <= 16'hC369;
11'h27C: o <= 16'hC356;
11'h27D: o <= 16'hC343;
11'h27E: o <= 16'hC331;
11'h27F: o <= 16'hC31E;
11'h280: o <= 16'hC30C;
11'h281: o <= 16'hC2F9;
11'h282: o <= 16'hC2E7;
11'h283: o <= 16'hC2D4;
11'h284: o <= 16'hC2C1;
11'h285: o <= 16'hC2AF;
11'h286: o <= 16'hC29C;
11'h287: o <= 16'hC28A;
11'h288: o <= 16'hC278;
11'h289: o <= 16'hC265;
11'h28A: o <= 16'hC253;
11'h28B: o <= 16'hC240;
11'h28C: o <= 16'hC22E;
11'h28D: o <= 16'hC21B;
11'h28E: o <= 16'hC209;
11'h28F: o <= 16'hC1F7;
11'h290: o <= 16'hC1E4;
11'h291: o <= 16'hC1D2;
11'h292: o <= 16'hC1C0;
11'h293: o <= 16'hC1AD;
11'h294: o <= 16'hC19B;
11'h295: o <= 16'hC189;
11'h296: o <= 16'hC176;
11'h297: o <= 16'hC164;
11'h298: o <= 16'hC152;
11'h299: o <= 16'hC140;
11'h29A: o <= 16'hC12D;
11'h29B: o <= 16'hC11B;
11'h29C: o <= 16'hC109;
11'h29D: o <= 16'hC0F7;
11'h29E: o <= 16'hC0E5;
11'h29F: o <= 16'hC0D2;
11'h2A0: o <= 16'hC0C0;
11'h2A1: o <= 16'hC0AE;
11'h2A2: o <= 16'hC09C;
11'h2A3: o <= 16'hC08A;
11'h2A4: o <= 16'hC078;
11'h2A5: o <= 16'hC066;
11'h2A6: o <= 16'hC054;
11'h2A7: o <= 16'hC042;
11'h2A8: o <= 16'hC030;
11'h2A9: o <= 16'hC01E;
11'h2AA: o <= 16'hC00C;
11'h2AB: o <= 16'hBFFA;
11'h2AC: o <= 16'hBFE8;
11'h2AD: o <= 16'hBFD6;
11'h2AE: o <= 16'hBFC4;
11'h2AF: o <= 16'hBFB2;
11'h2B0: o <= 16'hBFA0;
11'h2B1: o <= 16'hBF8E;
11'h2B2: o <= 16'hBF7C;
11'h2B3: o <= 16'hBF6A;
11'h2B4: o <= 16'hBF58;
11'h2B5: o <= 16'hBF46;
11'h2B6: o <= 16'hBF34;
11'h2B7: o <= 16'hBF22;
11'h2B8: o <= 16'hBF11;
11'h2B9: o <= 16'hBEFF;
11'h2BA: o <= 16'hBEED;
11'h2BB: o <= 16'hBEDB;
11'h2BC: o <= 16'hBEC9;
11'h2BD: o <= 16'hBEB8;
11'h2BE: o <= 16'hBEA6;
11'h2BF: o <= 16'hBE94;
11'h2C0: o <= 16'hBE82;
11'h2C1: o <= 16'hBE71;
11'h2C2: o <= 16'hBE5F;
11'h2C3: o <= 16'hBE4D;
11'h2C4: o <= 16'hBE3C;
11'h2C5: o <= 16'hBE2A;
11'h2C6: o <= 16'hBE18;
11'h2C7: o <= 16'hBE07;
11'h2C8: o <= 16'hBDF5;
11'h2C9: o <= 16'hBDE3;
11'h2CA: o <= 16'hBDD2;
11'h2CB: o <= 16'hBDC0;
11'h2CC: o <= 16'hBDAF;
11'h2CD: o <= 16'hBD9D;
11'h2CE: o <= 16'hBD8C;
11'h2CF: o <= 16'hBD7A;
11'h2D0: o <= 16'hBD69;
11'h2D1: o <= 16'hBD57;
11'h2D2: o <= 16'hBD46;
11'h2D3: o <= 16'hBD34;
11'h2D4: o <= 16'hBD23;
11'h2D5: o <= 16'hBD11;
11'h2D6: o <= 16'hBD00;
11'h2D7: o <= 16'hBCEE;
11'h2D8: o <= 16'hBCDD;
11'h2D9: o <= 16'hBCCB;
11'h2DA: o <= 16'hBCBA;
11'h2DB: o <= 16'hBCA9;
11'h2DC: o <= 16'hBC97;
11'h2DD: o <= 16'hBC86;
11'h2DE: o <= 16'hBC75;
11'h2DF: o <= 16'hBC63;
11'h2E0: o <= 16'hBC52;
11'h2E1: o <= 16'hBC41;
11'h2E2: o <= 16'hBC2F;
11'h2E3: o <= 16'hBC1E;
11'h2E4: o <= 16'hBC0D;
11'h2E5: o <= 16'hBBFB;
11'h2E6: o <= 16'hBBEA;
11'h2E7: o <= 16'hBBD9;
11'h2E8: o <= 16'hBBC8;
11'h2E9: o <= 16'hBBB7;
11'h2EA: o <= 16'hBBA5;
11'h2EB: o <= 16'hBB94;
11'h2EC: o <= 16'hBB83;
11'h2ED: o <= 16'hBB72;
11'h2EE: o <= 16'hBB61;
11'h2EF: o <= 16'hBB50;
11'h2F0: o <= 16'hBB3E;
11'h2F1: o <= 16'hBB2D;
11'h2F2: o <= 16'hBB1C;
11'h2F3: o <= 16'hBB0B;
11'h2F4: o <= 16'hBAFA;
11'h2F5: o <= 16'hBAE9;
11'h2F6: o <= 16'hBAD8;
11'h2F7: o <= 16'hBAC7;
11'h2F8: o <= 16'hBAB6;
11'h2F9: o <= 16'hBAA5;
11'h2FA: o <= 16'hBA94;
11'h2FB: o <= 16'hBA83;
11'h2FC: o <= 16'hBA72;
11'h2FD: o <= 16'hBA61;
11'h2FE: o <= 16'hBA50;
11'h2FF: o <= 16'hBA3F;
11'h300: o <= 16'hBA2E;
11'h301: o <= 16'hBA1D;
11'h302: o <= 16'hBA0C;
11'h303: o <= 16'hB9FB;
11'h304: o <= 16'hB9EA;
11'h305: o <= 16'hB9DA;
11'h306: o <= 16'hB9C9;
11'h307: o <= 16'hB9B8;
11'h308: o <= 16'hB9A7;
11'h309: o <= 16'hB996;
11'h30A: o <= 16'hB985;
11'h30B: o <= 16'hB975;
11'h30C: o <= 16'hB964;
11'h30D: o <= 16'hB953;
11'h30E: o <= 16'hB942;
11'h30F: o <= 16'hB932;
11'h310: o <= 16'hB921;
11'h311: o <= 16'hB910;
11'h312: o <= 16'hB8FF;
11'h313: o <= 16'hB8EF;
11'h314: o <= 16'hB8DE;
11'h315: o <= 16'hB8CD;
11'h316: o <= 16'hB8BD;
11'h317: o <= 16'hB8AC;
11'h318: o <= 16'hB89B;
11'h319: o <= 16'hB88B;
11'h31A: o <= 16'hB87A;
11'h31B: o <= 16'hB869;
11'h31C: o <= 16'hB859;
11'h31D: o <= 16'hB848;
11'h31E: o <= 16'hB838;
11'h31F: o <= 16'hB827;
11'h320: o <= 16'hB817;
11'h321: o <= 16'hB806;
11'h322: o <= 16'hB7F5;
11'h323: o <= 16'hB7E5;
11'h324: o <= 16'hB7D4;
11'h325: o <= 16'hB7C4;
11'h326: o <= 16'hB7B3;
11'h327: o <= 16'hB7A3;
11'h328: o <= 16'hB793;
11'h329: o <= 16'hB782;
11'h32A: o <= 16'hB772;
11'h32B: o <= 16'hB761;
11'h32C: o <= 16'hB751;
11'h32D: o <= 16'hB740;
11'h32E: o <= 16'hB730;
11'h32F: o <= 16'hB720;
11'h330: o <= 16'hB70F;
11'h331: o <= 16'hB6FF;
11'h332: o <= 16'hB6EF;
11'h333: o <= 16'hB6DE;
11'h334: o <= 16'hB6CE;
11'h335: o <= 16'hB6BE;
11'h336: o <= 16'hB6AD;
11'h337: o <= 16'hB69D;
11'h338: o <= 16'hB68D;
11'h339: o <= 16'hB67C;
11'h33A: o <= 16'hB66C;
11'h33B: o <= 16'hB65C;
11'h33C: o <= 16'hB64C;
11'h33D: o <= 16'hB63B;
11'h33E: o <= 16'hB62B;
11'h33F: o <= 16'hB61B;
11'h340: o <= 16'hB60B;
11'h341: o <= 16'hB5FB;
11'h342: o <= 16'hB5EB;
11'h343: o <= 16'hB5DA;
11'h344: o <= 16'hB5CA;
11'h345: o <= 16'hB5BA;
11'h346: o <= 16'hB5AA;
11'h347: o <= 16'hB59A;
11'h348: o <= 16'hB58A;
11'h349: o <= 16'hB57A;
11'h34A: o <= 16'hB56A;
11'h34B: o <= 16'hB55A;
11'h34C: o <= 16'hB54A;
11'h34D: o <= 16'hB539;
11'h34E: o <= 16'hB529;
11'h34F: o <= 16'hB519;
11'h350: o <= 16'hB509;
11'h351: o <= 16'hB4F9;
11'h352: o <= 16'hB4E9;
11'h353: o <= 16'hB4D9;
11'h354: o <= 16'hB4C9;
11'h355: o <= 16'hB4BA;
11'h356: o <= 16'hB4AA;
11'h357: o <= 16'hB49A;
11'h358: o <= 16'hB48A;
11'h359: o <= 16'hB47A;
11'h35A: o <= 16'hB46A;
11'h35B: o <= 16'hB45A;
11'h35C: o <= 16'hB44A;
11'h35D: o <= 16'hB43A;
11'h35E: o <= 16'hB42A;
11'h35F: o <= 16'hB41B;
11'h360: o <= 16'hB40B;
11'h361: o <= 16'hB3FB;
11'h362: o <= 16'hB3EB;
11'h363: o <= 16'hB3DB;
11'h364: o <= 16'hB3CC;
11'h365: o <= 16'hB3BC;
11'h366: o <= 16'hB3AC;
11'h367: o <= 16'hB39C;
11'h368: o <= 16'hB38C;
11'h369: o <= 16'hB37D;
11'h36A: o <= 16'hB36D;
11'h36B: o <= 16'hB35D;
11'h36C: o <= 16'hB34E;
11'h36D: o <= 16'hB33E;
11'h36E: o <= 16'hB32E;
11'h36F: o <= 16'hB31F;
11'h370: o <= 16'hB30F;
11'h371: o <= 16'hB2FF;
11'h372: o <= 16'hB2F0;
11'h373: o <= 16'hB2E0;
11'h374: o <= 16'hB2D0;
11'h375: o <= 16'hB2C1;
11'h376: o <= 16'hB2B1;
11'h377: o <= 16'hB2A2;
11'h378: o <= 16'hB292;
11'h379: o <= 16'hB282;
11'h37A: o <= 16'hB273;
11'h37B: o <= 16'hB263;
11'h37C: o <= 16'hB254;
11'h37D: o <= 16'hB244;
11'h37E: o <= 16'hB235;
11'h37F: o <= 16'hB225;
11'h380: o <= 16'hB216;
11'h381: o <= 16'hB206;
11'h382: o <= 16'hB1F7;
11'h383: o <= 16'hB1E7;
11'h384: o <= 16'hB1D8;
11'h385: o <= 16'hB1C8;
11'h386: o <= 16'hB1B9;
11'h387: o <= 16'hB1AA;
11'h388: o <= 16'hB19A;
11'h389: o <= 16'hB18B;
11'h38A: o <= 16'hB17B;
11'h38B: o <= 16'hB16C;
11'h38C: o <= 16'hB15D;
11'h38D: o <= 16'hB14D;
11'h38E: o <= 16'hB13E;
11'h38F: o <= 16'hB12F;
11'h390: o <= 16'hB11F;
11'h391: o <= 16'hB110;
11'h392: o <= 16'hB101;
11'h393: o <= 16'hB0F1;
11'h394: o <= 16'hB0E2;
11'h395: o <= 16'hB0D3;
11'h396: o <= 16'hB0C4;
11'h397: o <= 16'hB0B4;
11'h398: o <= 16'hB0A5;
11'h399: o <= 16'hB096;
11'h39A: o <= 16'hB087;
11'h39B: o <= 16'hB077;
11'h39C: o <= 16'hB068;
11'h39D: o <= 16'hB059;
11'h39E: o <= 16'hB04A;
11'h39F: o <= 16'hB03B;
11'h3A0: o <= 16'hB02C;
11'h3A1: o <= 16'hB01C;
11'h3A2: o <= 16'hB00D;
11'h3A3: o <= 16'hAFFE;
11'h3A4: o <= 16'hAFEF;
11'h3A5: o <= 16'hAFE0;
11'h3A6: o <= 16'hAFD1;
11'h3A7: o <= 16'hAFC2;
11'h3A8: o <= 16'hAFB3;
11'h3A9: o <= 16'hAFA4;
11'h3AA: o <= 16'hAF95;
11'h3AB: o <= 16'hAF85;
11'h3AC: o <= 16'hAF76;
11'h3AD: o <= 16'hAF67;
11'h3AE: o <= 16'hAF58;
11'h3AF: o <= 16'hAF49;
11'h3B0: o <= 16'hAF3A;
11'h3B1: o <= 16'hAF2B;
11'h3B2: o <= 16'hAF1C;
11'h3B3: o <= 16'hAF0D;
11'h3B4: o <= 16'hAEFE;
11'h3B5: o <= 16'hAEF0;
11'h3B6: o <= 16'hAEE1;
11'h3B7: o <= 16'hAED2;
11'h3B8: o <= 16'hAEC3;
11'h3B9: o <= 16'hAEB4;
11'h3BA: o <= 16'hAEA5;
11'h3BB: o <= 16'hAE96;
11'h3BC: o <= 16'hAE87;
11'h3BD: o <= 16'hAE78;
11'h3BE: o <= 16'hAE69;
11'h3BF: o <= 16'hAE5B;
11'h3C0: o <= 16'hAE4C;
11'h3C1: o <= 16'hAE3D;
11'h3C2: o <= 16'hAE2E;
11'h3C3: o <= 16'hAE1F;
11'h3C4: o <= 16'hAE10;
11'h3C5: o <= 16'hAE02;
11'h3C6: o <= 16'hADF3;
11'h3C7: o <= 16'hADE4;
11'h3C8: o <= 16'hADD5;
11'h3C9: o <= 16'hADC7;
11'h3CA: o <= 16'hADB8;
11'h3CB: o <= 16'hADA9;
11'h3CC: o <= 16'hAD9A;
11'h3CD: o <= 16'hAD8C;
11'h3CE: o <= 16'hAD7D;
11'h3CF: o <= 16'hAD6E;
11'h3D0: o <= 16'hAD60;
11'h3D1: o <= 16'hAD51;
11'h3D2: o <= 16'hAD42;
11'h3D3: o <= 16'hAD34;
11'h3D4: o <= 16'hAD25;
11'h3D5: o <= 16'hAD16;
11'h3D6: o <= 16'hAD08;
11'h3D7: o <= 16'hACF9;
11'h3D8: o <= 16'hACEB;
11'h3D9: o <= 16'hACDC;
11'h3DA: o <= 16'hACCD;
11'h3DB: o <= 16'hACBF;
11'h3DC: o <= 16'hACB0;
11'h3DD: o <= 16'hACA2;
11'h3DE: o <= 16'hAC93;
11'h3DF: o <= 16'hAC85;
11'h3E0: o <= 16'hAC76;
11'h3E1: o <= 16'hAC68;
11'h3E2: o <= 16'hAC59;
11'h3E3: o <= 16'hAC4B;
11'h3E4: o <= 16'hAC3C;
11'h3E5: o <= 16'hAC2E;
11'h3E6: o <= 16'hAC1F;
11'h3E7: o <= 16'hAC11;
11'h3E8: o <= 16'hAC02;
11'h3E9: o <= 16'hABF4;
11'h3EA: o <= 16'hABE5;
11'h3EB: o <= 16'hABD7;
11'h3EC: o <= 16'hABC8;
11'h3ED: o <= 16'hABBA;
11'h3EE: o <= 16'hABAC;
11'h3EF: o <= 16'hAB9D;
11'h3F0: o <= 16'hAB8F;
11'h3F1: o <= 16'hAB81;
11'h3F2: o <= 16'hAB72;
11'h3F3: o <= 16'hAB64;
11'h3F4: o <= 16'hAB56;
11'h3F5: o <= 16'hAB47;
11'h3F6: o <= 16'hAB39;
11'h3F7: o <= 16'hAB2B;
11'h3F8: o <= 16'hAB1C;
11'h3F9: o <= 16'hAB0E;
11'h3FA: o <= 16'hAB00;
11'h3FB: o <= 16'hAAF1;
11'h3FC: o <= 16'hAAE3;
11'h3FD: o <= 16'hAAD5;
11'h3FE: o <= 16'hAAC7;
11'h3FF: o <= 16'hAAB8;
11'h400: o <= 16'hAAAA;
11'h401: o <= 16'hAA9C;
11'h402: o <= 16'hAA8E;
11'h403: o <= 16'hAA80;
11'h404: o <= 16'hAA71;
11'h405: o <= 16'hAA63;
11'h406: o <= 16'hAA55;
11'h407: o <= 16'hAA47;
11'h408: o <= 16'hAA39;
11'h409: o <= 16'hAA2B;
11'h40A: o <= 16'hAA1C;
11'h40B: o <= 16'hAA0E;
11'h40C: o <= 16'hAA00;
11'h40D: o <= 16'hA9F2;
11'h40E: o <= 16'hA9E4;
11'h40F: o <= 16'hA9D6;
11'h410: o <= 16'hA9C8;
11'h411: o <= 16'hA9BA;
11'h412: o <= 16'hA9AC;
11'h413: o <= 16'hA99E;
11'h414: o <= 16'hA990;
11'h415: o <= 16'hA982;
11'h416: o <= 16'hA974;
11'h417: o <= 16'hA965;
11'h418: o <= 16'hA957;
11'h419: o <= 16'hA949;
11'h41A: o <= 16'hA93B;
11'h41B: o <= 16'hA92E;
11'h41C: o <= 16'hA920;
11'h41D: o <= 16'hA912;
11'h41E: o <= 16'hA904;
11'h41F: o <= 16'hA8F6;
11'h420: o <= 16'hA8E8;
11'h421: o <= 16'hA8DA;
11'h422: o <= 16'hA8CC;
11'h423: o <= 16'hA8BE;
11'h424: o <= 16'hA8B0;
11'h425: o <= 16'hA8A2;
11'h426: o <= 16'hA894;
11'h427: o <= 16'hA886;
11'h428: o <= 16'hA879;
11'h429: o <= 16'hA86B;
11'h42A: o <= 16'hA85D;
11'h42B: o <= 16'hA84F;
11'h42C: o <= 16'hA841;
11'h42D: o <= 16'hA833;
11'h42E: o <= 16'hA826;
11'h42F: o <= 16'hA818;
11'h430: o <= 16'hA80A;
11'h431: o <= 16'hA7FC;
11'h432: o <= 16'hA7EE;
11'h433: o <= 16'hA7E1;
11'h434: o <= 16'hA7D3;
11'h435: o <= 16'hA7C5;
11'h436: o <= 16'hA7B7;
11'h437: o <= 16'hA7AA;
11'h438: o <= 16'hA79C;
11'h439: o <= 16'hA78E;
11'h43A: o <= 16'hA781;
11'h43B: o <= 16'hA773;
11'h43C: o <= 16'hA765;
11'h43D: o <= 16'hA758;
11'h43E: o <= 16'hA74A;
11'h43F: o <= 16'hA73C;
11'h440: o <= 16'hA72F;
11'h441: o <= 16'hA721;
11'h442: o <= 16'hA713;
11'h443: o <= 16'hA706;
11'h444: o <= 16'hA6F8;
11'h445: o <= 16'hA6EA;
11'h446: o <= 16'hA6DD;
11'h447: o <= 16'hA6CF;
11'h448: o <= 16'hA6C2;
11'h449: o <= 16'hA6B4;
11'h44A: o <= 16'hA6A6;
11'h44B: o <= 16'hA699;
11'h44C: o <= 16'hA68B;
11'h44D: o <= 16'hA67E;
11'h44E: o <= 16'hA670;
11'h44F: o <= 16'hA663;
11'h450: o <= 16'hA655;
11'h451: o <= 16'hA648;
11'h452: o <= 16'hA63A;
11'h453: o <= 16'hA62D;
11'h454: o <= 16'hA61F;
11'h455: o <= 16'hA612;
11'h456: o <= 16'hA604;
11'h457: o <= 16'hA5F7;
11'h458: o <= 16'hA5E9;
11'h459: o <= 16'hA5DC;
11'h45A: o <= 16'hA5CF;
11'h45B: o <= 16'hA5C1;
11'h45C: o <= 16'hA5B4;
11'h45D: o <= 16'hA5A6;
11'h45E: o <= 16'hA599;
11'h45F: o <= 16'hA58C;
11'h460: o <= 16'hA57E;
11'h461: o <= 16'hA571;
11'h462: o <= 16'hA563;
11'h463: o <= 16'hA556;
11'h464: o <= 16'hA549;
11'h465: o <= 16'hA53B;
11'h466: o <= 16'hA52E;
11'h467: o <= 16'hA521;
11'h468: o <= 16'hA513;
11'h469: o <= 16'hA506;
11'h46A: o <= 16'hA4F9;
11'h46B: o <= 16'hA4EC;
11'h46C: o <= 16'hA4DE;
11'h46D: o <= 16'hA4D1;
11'h46E: o <= 16'hA4C4;
11'h46F: o <= 16'hA4B7;
11'h470: o <= 16'hA4A9;
11'h471: o <= 16'hA49C;
11'h472: o <= 16'hA48F;
11'h473: o <= 16'hA482;
11'h474: o <= 16'hA474;
11'h475: o <= 16'hA467;
11'h476: o <= 16'hA45A;
11'h477: o <= 16'hA44D;
11'h478: o <= 16'hA440;
11'h479: o <= 16'hA432;
11'h47A: o <= 16'hA425;
11'h47B: o <= 16'hA418;
11'h47C: o <= 16'hA40B;
11'h47D: o <= 16'hA3FE;
11'h47E: o <= 16'hA3F1;
11'h47F: o <= 16'hA3E4;
11'h480: o <= 16'hA3D7;
11'h481: o <= 16'hA3C9;
11'h482: o <= 16'hA3BC;
11'h483: o <= 16'hA3AF;
11'h484: o <= 16'hA3A2;
11'h485: o <= 16'hA395;
11'h486: o <= 16'hA388;
11'h487: o <= 16'hA37B;
11'h488: o <= 16'hA36E;
11'h489: o <= 16'hA361;
11'h48A: o <= 16'hA354;
11'h48B: o <= 16'hA347;
11'h48C: o <= 16'hA33A;
11'h48D: o <= 16'hA32D;
11'h48E: o <= 16'hA320;
11'h48F: o <= 16'hA313;
11'h490: o <= 16'hA306;
11'h491: o <= 16'hA2F9;
11'h492: o <= 16'hA2EC;
11'h493: o <= 16'hA2DF;
11'h494: o <= 16'hA2D2;
11'h495: o <= 16'hA2C5;
11'h496: o <= 16'hA2B8;
11'h497: o <= 16'hA2AB;
11'h498: o <= 16'hA29E;
11'h499: o <= 16'hA291;
11'h49A: o <= 16'hA284;
11'h49B: o <= 16'hA278;
11'h49C: o <= 16'hA26B;
11'h49D: o <= 16'hA25E;
11'h49E: o <= 16'hA251;
11'h49F: o <= 16'hA244;
11'h4A0: o <= 16'hA237;
11'h4A1: o <= 16'hA22A;
11'h4A2: o <= 16'hA21E;
11'h4A3: o <= 16'hA211;
11'h4A4: o <= 16'hA204;
11'h4A5: o <= 16'hA1F7;
11'h4A6: o <= 16'hA1EA;
11'h4A7: o <= 16'hA1DE;
11'h4A8: o <= 16'hA1D1;
11'h4A9: o <= 16'hA1C4;
11'h4AA: o <= 16'hA1B7;
11'h4AB: o <= 16'hA1AA;
11'h4AC: o <= 16'hA19E;
11'h4AD: o <= 16'hA191;
11'h4AE: o <= 16'hA184;
11'h4AF: o <= 16'hA177;
11'h4B0: o <= 16'hA16B;
11'h4B1: o <= 16'hA15E;
11'h4B2: o <= 16'hA151;
11'h4B3: o <= 16'hA145;
11'h4B4: o <= 16'hA138;
11'h4B5: o <= 16'hA12B;
11'h4B6: o <= 16'hA11E;
11'h4B7: o <= 16'hA112;
11'h4B8: o <= 16'hA105;
11'h4B9: o <= 16'hA0F9;
11'h4BA: o <= 16'hA0EC;
11'h4BB: o <= 16'hA0DF;
11'h4BC: o <= 16'hA0D3;
11'h4BD: o <= 16'hA0C6;
11'h4BE: o <= 16'hA0B9;
11'h4BF: o <= 16'hA0AD;
11'h4C0: o <= 16'hA0A0;
11'h4C1: o <= 16'hA094;
11'h4C2: o <= 16'hA087;
11'h4C3: o <= 16'hA07A;
11'h4C4: o <= 16'hA06E;
11'h4C5: o <= 16'hA061;
11'h4C6: o <= 16'hA055;
11'h4C7: o <= 16'hA048;
11'h4C8: o <= 16'hA03C;
11'h4C9: o <= 16'hA02F;
11'h4CA: o <= 16'hA023;
11'h4CB: o <= 16'hA016;
11'h4CC: o <= 16'hA00A;
11'h4CD: o <= 16'h9FFD;
11'h4CE: o <= 16'h9FF1;
11'h4CF: o <= 16'h9FE4;
11'h4D0: o <= 16'h9FD8;
11'h4D1: o <= 16'h9FCB;
11'h4D2: o <= 16'h9FBF;
11'h4D3: o <= 16'h9FB2;
11'h4D4: o <= 16'h9FA6;
11'h4D5: o <= 16'h9F99;
11'h4D6: o <= 16'h9F8D;
11'h4D7: o <= 16'h9F80;
11'h4D8: o <= 16'h9F74;
11'h4D9: o <= 16'h9F68;
11'h4DA: o <= 16'h9F5B;
11'h4DB: o <= 16'h9F4F;
11'h4DC: o <= 16'h9F42;
11'h4DD: o <= 16'h9F36;
11'h4DE: o <= 16'h9F2A;
11'h4DF: o <= 16'h9F1D;
11'h4E0: o <= 16'h9F11;
11'h4E1: o <= 16'h9F05;
11'h4E2: o <= 16'h9EF8;
11'h4E3: o <= 16'h9EEC;
11'h4E4: o <= 16'h9EE0;
11'h4E5: o <= 16'h9ED3;
11'h4E6: o <= 16'h9EC7;
11'h4E7: o <= 16'h9EBB;
11'h4E8: o <= 16'h9EAE;
11'h4E9: o <= 16'h9EA2;
11'h4EA: o <= 16'h9E96;
11'h4EB: o <= 16'h9E89;
11'h4EC: o <= 16'h9E7D;
11'h4ED: o <= 16'h9E71;
11'h4EE: o <= 16'h9E65;
11'h4EF: o <= 16'h9E58;
11'h4F0: o <= 16'h9E4C;
11'h4F1: o <= 16'h9E40;
11'h4F2: o <= 16'h9E34;
11'h4F3: o <= 16'h9E28;
11'h4F4: o <= 16'h9E1B;
11'h4F5: o <= 16'h9E0F;
11'h4F6: o <= 16'h9E03;
11'h4F7: o <= 16'h9DF7;
11'h4F8: o <= 16'h9DEB;
11'h4F9: o <= 16'h9DDE;
11'h4FA: o <= 16'h9DD2;
11'h4FB: o <= 16'h9DC6;
11'h4FC: o <= 16'h9DBA;
11'h4FD: o <= 16'h9DAE;
11'h4FE: o <= 16'h9DA2;
11'h4FF: o <= 16'h9D95;
11'h500: o <= 16'h9D89;
11'h501: o <= 16'h9D7D;
11'h502: o <= 16'h9D71;
11'h503: o <= 16'h9D65;
11'h504: o <= 16'h9D59;
11'h505: o <= 16'h9D4D;
11'h506: o <= 16'h9D41;
11'h507: o <= 16'h9D35;
11'h508: o <= 16'h9D29;
11'h509: o <= 16'h9D1D;
11'h50A: o <= 16'h9D11;
11'h50B: o <= 16'h9D04;
11'h50C: o <= 16'h9CF8;
11'h50D: o <= 16'h9CEC;
11'h50E: o <= 16'h9CE0;
11'h50F: o <= 16'h9CD4;
11'h510: o <= 16'h9CC8;
11'h511: o <= 16'h9CBC;
11'h512: o <= 16'h9CB0;
11'h513: o <= 16'h9CA4;
11'h514: o <= 16'h9C98;
11'h515: o <= 16'h9C8C;
11'h516: o <= 16'h9C80;
11'h517: o <= 16'h9C75;
11'h518: o <= 16'h9C69;
11'h519: o <= 16'h9C5D;
11'h51A: o <= 16'h9C51;
11'h51B: o <= 16'h9C45;
11'h51C: o <= 16'h9C39;
11'h51D: o <= 16'h9C2D;
11'h51E: o <= 16'h9C21;
11'h51F: o <= 16'h9C15;
11'h520: o <= 16'h9C09;
11'h521: o <= 16'h9BFD;
11'h522: o <= 16'h9BF1;
11'h523: o <= 16'h9BE6;
11'h524: o <= 16'h9BDA;
11'h525: o <= 16'h9BCE;
11'h526: o <= 16'h9BC2;
11'h527: o <= 16'h9BB6;
11'h528: o <= 16'h9BAA;
11'h529: o <= 16'h9B9F;
11'h52A: o <= 16'h9B93;
11'h52B: o <= 16'h9B87;
11'h52C: o <= 16'h9B7B;
11'h52D: o <= 16'h9B6F;
11'h52E: o <= 16'h9B64;
11'h52F: o <= 16'h9B58;
11'h530: o <= 16'h9B4C;
11'h531: o <= 16'h9B40;
11'h532: o <= 16'h9B34;
11'h533: o <= 16'h9B29;
11'h534: o <= 16'h9B1D;
11'h535: o <= 16'h9B11;
11'h536: o <= 16'h9B05;
11'h537: o <= 16'h9AFA;
11'h538: o <= 16'h9AEE;
11'h539: o <= 16'h9AE2;
11'h53A: o <= 16'h9AD7;
11'h53B: o <= 16'h9ACB;
11'h53C: o <= 16'h9ABF;
11'h53D: o <= 16'h9AB3;
11'h53E: o <= 16'h9AA8;
11'h53F: o <= 16'h9A9C;
11'h540: o <= 16'h9A90;
11'h541: o <= 16'h9A85;
11'h542: o <= 16'h9A79;
11'h543: o <= 16'h9A6D;
11'h544: o <= 16'h9A62;
11'h545: o <= 16'h9A56;
11'h546: o <= 16'h9A4B;
11'h547: o <= 16'h9A3F;
11'h548: o <= 16'h9A33;
11'h549: o <= 16'h9A28;
11'h54A: o <= 16'h9A1C;
11'h54B: o <= 16'h9A11;
11'h54C: o <= 16'h9A05;
11'h54D: o <= 16'h99F9;
11'h54E: o <= 16'h99EE;
11'h54F: o <= 16'h99E2;
11'h550: o <= 16'h99D7;
11'h551: o <= 16'h99CB;
11'h552: o <= 16'h99C0;
11'h553: o <= 16'h99B4;
11'h554: o <= 16'h99A8;
11'h555: o <= 16'h999D;
11'h556: o <= 16'h9991;
11'h557: o <= 16'h9986;
11'h558: o <= 16'h997A;
11'h559: o <= 16'h996F;
11'h55A: o <= 16'h9963;
11'h55B: o <= 16'h9958;
11'h55C: o <= 16'h994C;
11'h55D: o <= 16'h9941;
11'h55E: o <= 16'h9936;
11'h55F: o <= 16'h992A;
11'h560: o <= 16'h991F;
11'h561: o <= 16'h9913;
11'h562: o <= 16'h9908;
11'h563: o <= 16'h98FC;
11'h564: o <= 16'h98F1;
11'h565: o <= 16'h98E5;
11'h566: o <= 16'h98DA;
11'h567: o <= 16'h98CF;
11'h568: o <= 16'h98C3;
11'h569: o <= 16'h98B8;
11'h56A: o <= 16'h98AC;
11'h56B: o <= 16'h98A1;
11'h56C: o <= 16'h9896;
11'h56D: o <= 16'h988A;
11'h56E: o <= 16'h987F;
11'h56F: o <= 16'h9874;
11'h570: o <= 16'h9868;
11'h571: o <= 16'h985D;
11'h572: o <= 16'h9852;
11'h573: o <= 16'h9846;
11'h574: o <= 16'h983B;
11'h575: o <= 16'h9830;
11'h576: o <= 16'h9824;
11'h577: o <= 16'h9819;
11'h578: o <= 16'h980E;
11'h579: o <= 16'h9802;
11'h57A: o <= 16'h97F7;
11'h57B: o <= 16'h97EC;
11'h57C: o <= 16'h97E1;
11'h57D: o <= 16'h97D5;
11'h57E: o <= 16'h97CA;
11'h57F: o <= 16'h97BF;
11'h580: o <= 16'h97B4;
11'h581: o <= 16'h97A8;
11'h582: o <= 16'h979D;
11'h583: o <= 16'h9792;
11'h584: o <= 16'h9787;
11'h585: o <= 16'h977C;
11'h586: o <= 16'h9770;
11'h587: o <= 16'h9765;
11'h588: o <= 16'h975A;
11'h589: o <= 16'h974F;
11'h58A: o <= 16'h9744;
11'h58B: o <= 16'h9738;
11'h58C: o <= 16'h972D;
11'h58D: o <= 16'h9722;
11'h58E: o <= 16'h9717;
11'h58F: o <= 16'h970C;
11'h590: o <= 16'h9701;
11'h591: o <= 16'h96F6;
11'h592: o <= 16'h96EA;
11'h593: o <= 16'h96DF;
11'h594: o <= 16'h96D4;
11'h595: o <= 16'h96C9;
11'h596: o <= 16'h96BE;
11'h597: o <= 16'h96B3;
11'h598: o <= 16'h96A8;
11'h599: o <= 16'h969D;
11'h59A: o <= 16'h9692;
11'h59B: o <= 16'h9687;
11'h59C: o <= 16'h967C;
11'h59D: o <= 16'h9670;
11'h59E: o <= 16'h9665;
11'h59F: o <= 16'h965A;
11'h5A0: o <= 16'h964F;
11'h5A1: o <= 16'h9644;
11'h5A2: o <= 16'h9639;
11'h5A3: o <= 16'h962E;
11'h5A4: o <= 16'h9623;
11'h5A5: o <= 16'h9618;
11'h5A6: o <= 16'h960D;
11'h5A7: o <= 16'h9602;
11'h5A8: o <= 16'h95F7;
11'h5A9: o <= 16'h95EC;
11'h5AA: o <= 16'h95E1;
11'h5AB: o <= 16'h95D6;
11'h5AC: o <= 16'h95CB;
11'h5AD: o <= 16'h95C0;
11'h5AE: o <= 16'h95B6;
11'h5AF: o <= 16'h95AB;
11'h5B0: o <= 16'h95A0;
11'h5B1: o <= 16'h9595;
11'h5B2: o <= 16'h958A;
11'h5B3: o <= 16'h957F;
11'h5B4: o <= 16'h9574;
11'h5B5: o <= 16'h9569;
11'h5B6: o <= 16'h955E;
11'h5B7: o <= 16'h9553;
11'h5B8: o <= 16'h9548;
11'h5B9: o <= 16'h953E;
11'h5BA: o <= 16'h9533;
11'h5BB: o <= 16'h9528;
11'h5BC: o <= 16'h951D;
11'h5BD: o <= 16'h9512;
11'h5BE: o <= 16'h9507;
11'h5BF: o <= 16'h94FC;
11'h5C0: o <= 16'h94F2;
11'h5C1: o <= 16'h94E7;
11'h5C2: o <= 16'h94DC;
11'h5C3: o <= 16'h94D1;
11'h5C4: o <= 16'h94C6;
11'h5C5: o <= 16'h94BB;
11'h5C6: o <= 16'h94B1;
11'h5C7: o <= 16'h94A6;
11'h5C8: o <= 16'h949B;
11'h5C9: o <= 16'h9490;
11'h5CA: o <= 16'h9486;
11'h5CB: o <= 16'h947B;
11'h5CC: o <= 16'h9470;
11'h5CD: o <= 16'h9465;
11'h5CE: o <= 16'h945A;
11'h5CF: o <= 16'h9450;
11'h5D0: o <= 16'h9445;
11'h5D1: o <= 16'h943A;
11'h5D2: o <= 16'h9430;
11'h5D3: o <= 16'h9425;
11'h5D4: o <= 16'h941A;
11'h5D5: o <= 16'h940F;
11'h5D6: o <= 16'h9405;
11'h5D7: o <= 16'h93FA;
11'h5D8: o <= 16'h93EF;
11'h5D9: o <= 16'h93E5;
11'h5DA: o <= 16'h93DA;
11'h5DB: o <= 16'h93CF;
11'h5DC: o <= 16'h93C5;
11'h5DD: o <= 16'h93BA;
11'h5DE: o <= 16'h93AF;
11'h5DF: o <= 16'h93A5;
11'h5E0: o <= 16'h939A;
11'h5E1: o <= 16'h938F;
11'h5E2: o <= 16'h9385;
11'h5E3: o <= 16'h937A;
11'h5E4: o <= 16'h9370;
11'h5E5: o <= 16'h9365;
11'h5E6: o <= 16'h935A;
11'h5E7: o <= 16'h9350;
11'h5E8: o <= 16'h9345;
11'h5E9: o <= 16'h933B;
11'h5EA: o <= 16'h9330;
11'h5EB: o <= 16'h9325;
11'h5EC: o <= 16'h931B;
11'h5ED: o <= 16'h9310;
11'h5EE: o <= 16'h9306;
11'h5EF: o <= 16'h92FB;
11'h5F0: o <= 16'h92F1;
11'h5F1: o <= 16'h92E6;
11'h5F2: o <= 16'h92DC;
11'h5F3: o <= 16'h92D1;
11'h5F4: o <= 16'h92C6;
11'h5F5: o <= 16'h92BC;
11'h5F6: o <= 16'h92B1;
11'h5F7: o <= 16'h92A7;
11'h5F8: o <= 16'h929C;
11'h5F9: o <= 16'h9292;
11'h5FA: o <= 16'h9287;
11'h5FB: o <= 16'h927D;
11'h5FC: o <= 16'h9272;
11'h5FD: o <= 16'h9268;
11'h5FE: o <= 16'h925E;
11'h5FF: o <= 16'h9253;
11'h600: o <= 16'h9249;
11'h601: o <= 16'h923E;
11'h602: o <= 16'h9234;
11'h603: o <= 16'h9229;
11'h604: o <= 16'h921F;
11'h605: o <= 16'h9214;
11'h606: o <= 16'h920A;
11'h607: o <= 16'h9200;
11'h608: o <= 16'h91F5;
11'h609: o <= 16'h91EB;
11'h60A: o <= 16'h91E0;
11'h60B: o <= 16'h91D6;
11'h60C: o <= 16'h91CC;
11'h60D: o <= 16'h91C1;
11'h60E: o <= 16'h91B7;
11'h60F: o <= 16'h91AD;
11'h610: o <= 16'h91A2;
11'h611: o <= 16'h9198;
11'h612: o <= 16'h918E;
11'h613: o <= 16'h9183;
11'h614: o <= 16'h9179;
11'h615: o <= 16'h916E;
11'h616: o <= 16'h9164;
11'h617: o <= 16'h915A;
11'h618: o <= 16'h9150;
11'h619: o <= 16'h9145;
11'h61A: o <= 16'h913B;
11'h61B: o <= 16'h9131;
11'h61C: o <= 16'h9126;
11'h61D: o <= 16'h911C;
11'h61E: o <= 16'h9112;
11'h61F: o <= 16'h9108;
11'h620: o <= 16'h90FD;
11'h621: o <= 16'h90F3;
11'h622: o <= 16'h90E9;
11'h623: o <= 16'h90DE;
11'h624: o <= 16'h90D4;
11'h625: o <= 16'h90CA;
11'h626: o <= 16'h90C0;
11'h627: o <= 16'h90B6;
11'h628: o <= 16'h90AB;
11'h629: o <= 16'h90A1;
11'h62A: o <= 16'h9097;
11'h62B: o <= 16'h908D;
11'h62C: o <= 16'h9082;
11'h62D: o <= 16'h9078;
11'h62E: o <= 16'h906E;
11'h62F: o <= 16'h9064;
11'h630: o <= 16'h905A;
11'h631: o <= 16'h9050;
11'h632: o <= 16'h9045;
11'h633: o <= 16'h903B;
11'h634: o <= 16'h9031;
11'h635: o <= 16'h9027;
11'h636: o <= 16'h901D;
11'h637: o <= 16'h9013;
11'h638: o <= 16'h9009;
11'h639: o <= 16'h8FFE;
11'h63A: o <= 16'h8FF4;
11'h63B: o <= 16'h8FEA;
11'h63C: o <= 16'h8FE0;
11'h63D: o <= 16'h8FD6;
11'h63E: o <= 16'h8FCC;
11'h63F: o <= 16'h8FC2;
11'h640: o <= 16'h8FB8;
11'h641: o <= 16'h8FAE;
11'h642: o <= 16'h8FA3;
11'h643: o <= 16'h8F99;
11'h644: o <= 16'h8F8F;
11'h645: o <= 16'h8F85;
11'h646: o <= 16'h8F7B;
11'h647: o <= 16'h8F71;
11'h648: o <= 16'h8F67;
11'h649: o <= 16'h8F5D;
11'h64A: o <= 16'h8F53;
11'h64B: o <= 16'h8F49;
11'h64C: o <= 16'h8F3F;
11'h64D: o <= 16'h8F35;
11'h64E: o <= 16'h8F2B;
11'h64F: o <= 16'h8F21;
11'h650: o <= 16'h8F17;
11'h651: o <= 16'h8F0D;
11'h652: o <= 16'h8F03;
11'h653: o <= 16'h8EF9;
11'h654: o <= 16'h8EEF;
11'h655: o <= 16'h8EE5;
11'h656: o <= 16'h8EDB;
11'h657: o <= 16'h8ED1;
11'h658: o <= 16'h8EC7;
11'h659: o <= 16'h8EBD;
11'h65A: o <= 16'h8EB3;
11'h65B: o <= 16'h8EA9;
11'h65C: o <= 16'h8E9F;
11'h65D: o <= 16'h8E95;
11'h65E: o <= 16'h8E8C;
11'h65F: o <= 16'h8E82;
11'h660: o <= 16'h8E78;
11'h661: o <= 16'h8E6E;
11'h662: o <= 16'h8E64;
11'h663: o <= 16'h8E5A;
11'h664: o <= 16'h8E50;
11'h665: o <= 16'h8E46;
11'h666: o <= 16'h8E3C;
11'h667: o <= 16'h8E32;
11'h668: o <= 16'h8E29;
11'h669: o <= 16'h8E1F;
11'h66A: o <= 16'h8E15;
11'h66B: o <= 16'h8E0B;
11'h66C: o <= 16'h8E01;
11'h66D: o <= 16'h8DF7;
11'h66E: o <= 16'h8DED;
11'h66F: o <= 16'h8DE4;
11'h670: o <= 16'h8DDA;
11'h671: o <= 16'h8DD0;
11'h672: o <= 16'h8DC6;
11'h673: o <= 16'h8DBC;
11'h674: o <= 16'h8DB3;
11'h675: o <= 16'h8DA9;
11'h676: o <= 16'h8D9F;
11'h677: o <= 16'h8D95;
11'h678: o <= 16'h8D8B;
11'h679: o <= 16'h8D82;
11'h67A: o <= 16'h8D78;
11'h67B: o <= 16'h8D6E;
11'h67C: o <= 16'h8D64;
11'h67D: o <= 16'h8D5B;
11'h67E: o <= 16'h8D51;
11'h67F: o <= 16'h8D47;
11'h680: o <= 16'h8D3D;
11'h681: o <= 16'h8D34;
11'h682: o <= 16'h8D2A;
11'h683: o <= 16'h8D20;
11'h684: o <= 16'h8D16;
11'h685: o <= 16'h8D0D;
11'h686: o <= 16'h8D03;
11'h687: o <= 16'h8CF9;
11'h688: o <= 16'h8CF0;
11'h689: o <= 16'h8CE6;
11'h68A: o <= 16'h8CDC;
11'h68B: o <= 16'h8CD2;
11'h68C: o <= 16'h8CC9;
11'h68D: o <= 16'h8CBF;
11'h68E: o <= 16'h8CB5;
11'h68F: o <= 16'h8CAC;
11'h690: o <= 16'h8CA2;
11'h691: o <= 16'h8C98;
11'h692: o <= 16'h8C8F;
11'h693: o <= 16'h8C85;
11'h694: o <= 16'h8C7C;
11'h695: o <= 16'h8C72;
11'h696: o <= 16'h8C68;
11'h697: o <= 16'h8C5F;
11'h698: o <= 16'h8C55;
11'h699: o <= 16'h8C4B;
11'h69A: o <= 16'h8C42;
11'h69B: o <= 16'h8C38;
11'h69C: o <= 16'h8C2F;
11'h69D: o <= 16'h8C25;
11'h69E: o <= 16'h8C1B;
11'h69F: o <= 16'h8C12;
11'h6A0: o <= 16'h8C08;
11'h6A1: o <= 16'h8BFF;
11'h6A2: o <= 16'h8BF5;
11'h6A3: o <= 16'h8BEC;
11'h6A4: o <= 16'h8BE2;
11'h6A5: o <= 16'h8BD8;
11'h6A6: o <= 16'h8BCF;
11'h6A7: o <= 16'h8BC5;
11'h6A8: o <= 16'h8BBC;
11'h6A9: o <= 16'h8BB2;
11'h6AA: o <= 16'h8BA9;
11'h6AB: o <= 16'h8B9F;
11'h6AC: o <= 16'h8B96;
11'h6AD: o <= 16'h8B8C;
11'h6AE: o <= 16'h8B83;
11'h6AF: o <= 16'h8B79;
11'h6B0: o <= 16'h8B70;
11'h6B1: o <= 16'h8B66;
11'h6B2: o <= 16'h8B5D;
11'h6B3: o <= 16'h8B53;
11'h6B4: o <= 16'h8B4A;
11'h6B5: o <= 16'h8B40;
11'h6B6: o <= 16'h8B37;
11'h6B7: o <= 16'h8B2D;
11'h6B8: o <= 16'h8B24;
11'h6B9: o <= 16'h8B1A;
11'h6BA: o <= 16'h8B11;
11'h6BB: o <= 16'h8B08;
11'h6BC: o <= 16'h8AFE;
11'h6BD: o <= 16'h8AF5;
11'h6BE: o <= 16'h8AEB;
11'h6BF: o <= 16'h8AE2;
11'h6C0: o <= 16'h8AD8;
11'h6C1: o <= 16'h8ACF;
11'h6C2: o <= 16'h8AC6;
11'h6C3: o <= 16'h8ABC;
11'h6C4: o <= 16'h8AB3;
11'h6C5: o <= 16'h8AA9;
11'h6C6: o <= 16'h8AA0;
11'h6C7: o <= 16'h8A97;
11'h6C8: o <= 16'h8A8D;
11'h6C9: o <= 16'h8A84;
11'h6CA: o <= 16'h8A7B;
11'h6CB: o <= 16'h8A71;
11'h6CC: o <= 16'h8A68;
11'h6CD: o <= 16'h8A5E;
11'h6CE: o <= 16'h8A55;
11'h6CF: o <= 16'h8A4C;
11'h6D0: o <= 16'h8A42;
11'h6D1: o <= 16'h8A39;
11'h6D2: o <= 16'h8A30;
11'h6D3: o <= 16'h8A26;
11'h6D4: o <= 16'h8A1D;
11'h6D5: o <= 16'h8A14;
11'h6D6: o <= 16'h8A0B;
11'h6D7: o <= 16'h8A01;
11'h6D8: o <= 16'h89F8;
11'h6D9: o <= 16'h89EF;
11'h6DA: o <= 16'h89E5;
11'h6DB: o <= 16'h89DC;
11'h6DC: o <= 16'h89D3;
11'h6DD: o <= 16'h89CA;
11'h6DE: o <= 16'h89C0;
11'h6DF: o <= 16'h89B7;
11'h6E0: o <= 16'h89AE;
11'h6E1: o <= 16'h89A4;
11'h6E2: o <= 16'h899B;
11'h6E3: o <= 16'h8992;
11'h6E4: o <= 16'h8989;
11'h6E5: o <= 16'h8980;
11'h6E6: o <= 16'h8976;
11'h6E7: o <= 16'h896D;
11'h6E8: o <= 16'h8964;
11'h6E9: o <= 16'h895B;
11'h6EA: o <= 16'h8951;
11'h6EB: o <= 16'h8948;
11'h6EC: o <= 16'h893F;
11'h6ED: o <= 16'h8936;
11'h6EE: o <= 16'h892D;
11'h6EF: o <= 16'h8923;
11'h6F0: o <= 16'h891A;
11'h6F1: o <= 16'h8911;
11'h6F2: o <= 16'h8908;
11'h6F3: o <= 16'h88FF;
11'h6F4: o <= 16'h88F6;
11'h6F5: o <= 16'h88EC;
11'h6F6: o <= 16'h88E3;
11'h6F7: o <= 16'h88DA;
11'h6F8: o <= 16'h88D1;
11'h6F9: o <= 16'h88C8;
11'h6FA: o <= 16'h88BF;
11'h6FB: o <= 16'h88B6;
11'h6FC: o <= 16'h88AC;
11'h6FD: o <= 16'h88A3;
11'h6FE: o <= 16'h889A;
11'h6FF: o <= 16'h8891;
11'h700: o <= 16'h8888;
11'h701: o <= 16'h887F;
11'h702: o <= 16'h8876;
11'h703: o <= 16'h886D;
11'h704: o <= 16'h8864;
11'h705: o <= 16'h885B;
11'h706: o <= 16'h8852;
11'h707: o <= 16'h8848;
11'h708: o <= 16'h883F;
11'h709: o <= 16'h8836;
11'h70A: o <= 16'h882D;
11'h70B: o <= 16'h8824;
11'h70C: o <= 16'h881B;
11'h70D: o <= 16'h8812;
11'h70E: o <= 16'h8809;
11'h70F: o <= 16'h8800;
11'h710: o <= 16'h87F7;
11'h711: o <= 16'h87EE;
11'h712: o <= 16'h87E5;
11'h713: o <= 16'h87DC;
11'h714: o <= 16'h87D3;
11'h715: o <= 16'h87CA;
11'h716: o <= 16'h87C1;
11'h717: o <= 16'h87B8;
11'h718: o <= 16'h87AF;
11'h719: o <= 16'h87A6;
11'h71A: o <= 16'h879D;
11'h71B: o <= 16'h8794;
11'h71C: o <= 16'h878B;
11'h71D: o <= 16'h8782;
11'h71E: o <= 16'h8779;
11'h71F: o <= 16'h8770;
11'h720: o <= 16'h8767;
11'h721: o <= 16'h875E;
11'h722: o <= 16'h8755;
11'h723: o <= 16'h874C;
11'h724: o <= 16'h8743;
11'h725: o <= 16'h873A;
11'h726: o <= 16'h8732;
11'h727: o <= 16'h8729;
11'h728: o <= 16'h8720;
11'h729: o <= 16'h8717;
11'h72A: o <= 16'h870E;
11'h72B: o <= 16'h8705;
11'h72C: o <= 16'h86FC;
11'h72D: o <= 16'h86F3;
11'h72E: o <= 16'h86EA;
11'h72F: o <= 16'h86E1;
11'h730: o <= 16'h86D9;
11'h731: o <= 16'h86D0;
11'h732: o <= 16'h86C7;
11'h733: o <= 16'h86BE;
11'h734: o <= 16'h86B5;
11'h735: o <= 16'h86AC;
11'h736: o <= 16'h86A3;
11'h737: o <= 16'h869A;
11'h738: o <= 16'h8692;
11'h739: o <= 16'h8689;
11'h73A: o <= 16'h8680;
11'h73B: o <= 16'h8677;
11'h73C: o <= 16'h866E;
11'h73D: o <= 16'h8665;
11'h73E: o <= 16'h865D;
11'h73F: o <= 16'h8654;
11'h740: o <= 16'h864B;
11'h741: o <= 16'h8642;
11'h742: o <= 16'h8639;
11'h743: o <= 16'h8631;
11'h744: o <= 16'h8628;
11'h745: o <= 16'h861F;
11'h746: o <= 16'h8616;
11'h747: o <= 16'h860E;
11'h748: o <= 16'h8605;
11'h749: o <= 16'h85FC;
11'h74A: o <= 16'h85F3;
11'h74B: o <= 16'h85EA;
11'h74C: o <= 16'h85E2;
11'h74D: o <= 16'h85D9;
11'h74E: o <= 16'h85D0;
11'h74F: o <= 16'h85C7;
11'h750: o <= 16'h85BF;
11'h751: o <= 16'h85B6;
11'h752: o <= 16'h85AD;
11'h753: o <= 16'h85A5;
11'h754: o <= 16'h859C;
11'h755: o <= 16'h8593;
11'h756: o <= 16'h858A;
11'h757: o <= 16'h8582;
11'h758: o <= 16'h8579;
11'h759: o <= 16'h8570;
11'h75A: o <= 16'h8568;
11'h75B: o <= 16'h855F;
11'h75C: o <= 16'h8556;
11'h75D: o <= 16'h854E;
11'h75E: o <= 16'h8545;
11'h75F: o <= 16'h853C;
11'h760: o <= 16'h8534;
11'h761: o <= 16'h852B;
11'h762: o <= 16'h8522;
11'h763: o <= 16'h851A;
11'h764: o <= 16'h8511;
11'h765: o <= 16'h8508;
11'h766: o <= 16'h8500;
11'h767: o <= 16'h84F7;
11'h768: o <= 16'h84EE;
11'h769: o <= 16'h84E6;
11'h76A: o <= 16'h84DD;
11'h76B: o <= 16'h84D4;
11'h76C: o <= 16'h84CC;
11'h76D: o <= 16'h84C3;
11'h76E: o <= 16'h84BB;
11'h76F: o <= 16'h84B2;
11'h770: o <= 16'h84A9;
11'h771: o <= 16'h84A1;
11'h772: o <= 16'h8498;
11'h773: o <= 16'h8490;
11'h774: o <= 16'h8487;
11'h775: o <= 16'h847F;
11'h776: o <= 16'h8476;
11'h777: o <= 16'h846D;
11'h778: o <= 16'h8465;
11'h779: o <= 16'h845C;
11'h77A: o <= 16'h8454;
11'h77B: o <= 16'h844B;
11'h77C: o <= 16'h8443;
11'h77D: o <= 16'h843A;
11'h77E: o <= 16'h8432;
11'h77F: o <= 16'h8429;
11'h780: o <= 16'h8421;
11'h781: o <= 16'h8418;
11'h782: o <= 16'h840F;
11'h783: o <= 16'h8407;
11'h784: o <= 16'h83FE;
11'h785: o <= 16'h83F6;
11'h786: o <= 16'h83ED;
11'h787: o <= 16'h83E5;
11'h788: o <= 16'h83DC;
11'h789: o <= 16'h83D4;
11'h78A: o <= 16'h83CC;
11'h78B: o <= 16'h83C3;
11'h78C: o <= 16'h83BB;
11'h78D: o <= 16'h83B2;
11'h78E: o <= 16'h83AA;
11'h78F: o <= 16'h83A1;
11'h790: o <= 16'h8399;
11'h791: o <= 16'h8390;
11'h792: o <= 16'h8388;
11'h793: o <= 16'h837F;
11'h794: o <= 16'h8377;
11'h795: o <= 16'h836E;
11'h796: o <= 16'h8366;
11'h797: o <= 16'h835E;
11'h798: o <= 16'h8355;
11'h799: o <= 16'h834D;
11'h79A: o <= 16'h8344;
11'h79B: o <= 16'h833C;
11'h79C: o <= 16'h8334;
11'h79D: o <= 16'h832B;
11'h79E: o <= 16'h8323;
11'h79F: o <= 16'h831A;
11'h7A0: o <= 16'h8312;
11'h7A1: o <= 16'h830A;
11'h7A2: o <= 16'h8301;
11'h7A3: o <= 16'h82F9;
11'h7A4: o <= 16'h82F0;
11'h7A5: o <= 16'h82E8;
11'h7A6: o <= 16'h82E0;
11'h7A7: o <= 16'h82D7;
11'h7A8: o <= 16'h82CF;
11'h7A9: o <= 16'h82C7;
11'h7AA: o <= 16'h82BE;
11'h7AB: o <= 16'h82B6;
11'h7AC: o <= 16'h82AE;
11'h7AD: o <= 16'h82A5;
11'h7AE: o <= 16'h829D;
11'h7AF: o <= 16'h8295;
11'h7B0: o <= 16'h828C;
11'h7B1: o <= 16'h8284;
11'h7B2: o <= 16'h827C;
11'h7B3: o <= 16'h8273;
11'h7B4: o <= 16'h826B;
11'h7B5: o <= 16'h8263;
11'h7B6: o <= 16'h825A;
11'h7B7: o <= 16'h8252;
11'h7B8: o <= 16'h824A;
11'h7B9: o <= 16'h8242;
11'h7BA: o <= 16'h8239;
11'h7BB: o <= 16'h8231;
11'h7BC: o <= 16'h8229;
11'h7BD: o <= 16'h8220;
11'h7BE: o <= 16'h8218;
11'h7BF: o <= 16'h8210;
11'h7C0: o <= 16'h8208;
11'h7C1: o <= 16'h81FF;
11'h7C2: o <= 16'h81F7;
11'h7C3: o <= 16'h81EF;
11'h7C4: o <= 16'h81E7;
11'h7C5: o <= 16'h81DE;
11'h7C6: o <= 16'h81D6;
11'h7C7: o <= 16'h81CE;
11'h7C8: o <= 16'h81C6;
11'h7C9: o <= 16'h81BD;
11'h7CA: o <= 16'h81B5;
11'h7CB: o <= 16'h81AD;
11'h7CC: o <= 16'h81A5;
11'h7CD: o <= 16'h819D;
11'h7CE: o <= 16'h8194;
11'h7CF: o <= 16'h818C;
11'h7D0: o <= 16'h8184;
11'h7D1: o <= 16'h817C;
11'h7D2: o <= 16'h8174;
11'h7D3: o <= 16'h816B;
11'h7D4: o <= 16'h8163;
11'h7D5: o <= 16'h815B;
11'h7D6: o <= 16'h8153;
11'h7D7: o <= 16'h814B;
11'h7D8: o <= 16'h8143;
11'h7D9: o <= 16'h813A;
11'h7DA: o <= 16'h8132;
11'h7DB: o <= 16'h812A;
11'h7DC: o <= 16'h8122;
11'h7DD: o <= 16'h811A;
11'h7DE: o <= 16'h8112;
11'h7DF: o <= 16'h810A;
11'h7E0: o <= 16'h8102;
11'h7E1: o <= 16'h80F9;
11'h7E2: o <= 16'h80F1;
11'h7E3: o <= 16'h80E9;
11'h7E4: o <= 16'h80E1;
11'h7E5: o <= 16'h80D9;
11'h7E6: o <= 16'h80D1;
11'h7E7: o <= 16'h80C9;
11'h7E8: o <= 16'h80C1;
11'h7E9: o <= 16'h80B9;
11'h7EA: o <= 16'h80B0;
11'h7EB: o <= 16'h80A8;
11'h7EC: o <= 16'h80A0;
11'h7ED: o <= 16'h8098;
11'h7EE: o <= 16'h8090;
11'h7EF: o <= 16'h8088;
11'h7F0: o <= 16'h8080;
11'h7F1: o <= 16'h8078;
11'h7F2: o <= 16'h8070;
11'h7F3: o <= 16'h8068;
11'h7F4: o <= 16'h8060;
11'h7F5: o <= 16'h8058;
11'h7F6: o <= 16'h8050;
11'h7F7: o <= 16'h8048;
11'h7F8: o <= 16'h8040;
11'h7F9: o <= 16'h8038;
11'h7FA: o <= 16'h8030;
11'h7FB: o <= 16'h8028;
11'h7FC: o <= 16'h8020;
11'h7FD: o <= 16'h8018;
11'h7FE: o <= 16'h8010;
11'h7FF: o <= 16'h8008;
endcase
endmodule
