module rtf64ss();

endmodule
