module GridRouter();
endmodule
