// ============================================================================
//        __
//   \\__/ o\    (C) 2017-2019  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	fpRsqrte.v
//		- reciprocal square root estimate
//
//
// This source file is free software: you can redistribute it and/or modify 
// it under the terms of the GNU Lesser General Public License as published 
// by the Free Software Foundation, either version 3 of the License, or     
// (at your option) any later version.                                      
//                                                                          
// This source file is distributed in the hope that it will be useful,      
// but WITHOUT ANY WARRANTY; without even the implied warranty of           
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the            
// GNU General Public License for more details.                             
//                                                                          
// You should have received a copy of the GNU General Public License        
// along with this program.  If not, see <http://www.gnu.org/licenses/>.    
//
//
// ============================================================================

`include "fp_defines.v"

`define POINT5			32'h3F000000
`define ONEPOINT5		32'h3FC00000
`define FRSQRTE_MAGIC		32'h5f3759df

//`define RSQRT_SM		1'b1
`define RSQRT_TBL		1'b1

module fpRsqrte(clk, ce, ld, a, o);
parameter WID = 80;
`include "fpSize.sv"
input clk;
input ce;
input ld;
input [WID-1:0] a;
output reg [WID-1:0] o;

// An implementation of the approximation used in the Quake game.

wire [31:0] x2, x2yy, x2yy1p5;
wire [31:0] y, yy;
`ifdef RSQRT_TBL
// Reciprocal square root estimate using lookup table.

reg [15:0] RsqrteLUT2 [0:67];
reg [15:0] RsqrteLUT [0:8191];

initial begin
// This table stores the top 17 bits of the reciprocal square root estimate.
// (The sign bit is not stored).
// This table has two purposes. 1) The first 8129 entries of a 16k word lookup
// table are all infinity values, since they are the reciprocal of really
// small numbers. That means there's no real need to store those values in a
// lookup table. However that leaves about 64 "extra" values beyond what an
// 8192 entry lookup table could hold. So these values are stored in a smaller
// 68-entry lookup table. 2) A handful of values require the MSB of the
// exponent to be set. They won't fit in the 8192 entry table. Fortunately
// there are only four values like that.
// 
RsqrteLUT2[0] = 16'h7f84;
RsqrteLUT2[1] = 16'h7f88;
RsqrteLUT2[2] = 16'h7f8c;
RsqrteLUT2[3] = 16'h7f90;
RsqrteLUT2[4] = 16'h7f94;
RsqrteLUT2[5] = 16'h7f98;
RsqrteLUT2[6] = 16'h7f9c;
RsqrteLUT2[7] = 16'h7fa0;
RsqrteLUT2[8] = 16'h7fa4;
RsqrteLUT2[9] = 16'h7fa8;
RsqrteLUT2[10] = 16'h7fac;
RsqrteLUT2[11] = 16'h7fb0;
RsqrteLUT2[12] = 16'h7fb4;
RsqrteLUT2[13] = 16'h7fb8;
RsqrteLUT2[14] = 16'h7fbc;
RsqrteLUT2[15] = 16'h7fc0;
RsqrteLUT2[16] = 16'h7fc4;
RsqrteLUT2[17] = 16'h7fc8;
RsqrteLUT2[18] = 16'h7fcc;
RsqrteLUT2[19] = 16'h7fd0;
RsqrteLUT2[20] = 16'h7fd4;
RsqrteLUT2[21] = 16'h7fd8;
RsqrteLUT2[22] = 16'h7fdc;
RsqrteLUT2[23] = 16'h7fe0;
RsqrteLUT2[24] = 16'h7fe4;
RsqrteLUT2[25] = 16'h7fe8;
RsqrteLUT2[26] = 16'h7fec;
RsqrteLUT2[27] = 16'h7ff0;
RsqrteLUT2[28] = 16'h7ff4;
RsqrteLUT2[29] = 16'h7ff8;
RsqrteLUT2[30] = 16'h7ffc;
RsqrteLUT2[31] = 16'h7f80;
RsqrteLUT2[32] = 16'h7f84;
RsqrteLUT2[33] = 16'h7f88;
RsqrteLUT2[34] = 16'h7f8c;
RsqrteLUT2[35] = 16'h7f90;
RsqrteLUT2[36] = 16'h7f94;
RsqrteLUT2[37] = 16'h7f98;
RsqrteLUT2[38] = 16'h7f9c;
RsqrteLUT2[39] = 16'h7fa0;
RsqrteLUT2[40] = 16'h7fa4;
RsqrteLUT2[41] = 16'h7fa8;
RsqrteLUT2[42] = 16'h7fac;
RsqrteLUT2[43] = 16'h7fb0;
RsqrteLUT2[44] = 16'h7fb4;
RsqrteLUT2[45] = 16'h7fb8;
RsqrteLUT2[46] = 16'h7fbc;
RsqrteLUT2[47] = 16'h7fc0;
RsqrteLUT2[48] = 16'h7fc4;
RsqrteLUT2[49] = 16'h7fc8;
RsqrteLUT2[50] = 16'h7fcc;
RsqrteLUT2[51] = 16'h7fd0;
RsqrteLUT2[52] = 16'h7fd4;
RsqrteLUT2[53] = 16'h7fd8;
RsqrteLUT2[54] = 16'h7fdc;
RsqrteLUT2[55] = 16'h7fe0;
RsqrteLUT2[56] = 16'h7fe4;
RsqrteLUT2[57] = 16'h7fe8;
RsqrteLUT2[58] = 16'h7fec;
RsqrteLUT2[59] = 16'h7ff0;
RsqrteLUT2[60] = 16'h7ff4;
RsqrteLUT2[61] = 16'h7ff8;
RsqrteLUT2[62] = 16'h7ffc;
RsqrteLUT2[63] = 16'h7f00;
RsqrteLUT2[64] = 16'h8100;
RsqrteLUT2[65] = 16'h806a;
RsqrteLUT2[66] = 16'h8027;
RsqrteLUT2[67] = 16'h8000;
// This table stores the top 18 bits of the reciprocal square root estimate
// for 32-bit single precision values. The sign bit is not stored. Also the
// MSB of the exponent is not stored (for this table it's always zero). That
// allows the top 9 bits of the mantissa to be stored. The final result won't
// be accurate to more than six bits however, as that is the number of bits
// from the mantissa used to lookup the result.
RsqrteLUT[5] = 16'hff93;
RsqrteLUT[6] = 16'hff44;
RsqrteLUT[7] = 16'hff06;
RsqrteLUT[8] = 16'hfed4;
RsqrteLUT[9] = 16'hfeaa;
RsqrteLUT[10] = 16'hfe87;
RsqrteLUT[11] = 16'hfe69;
RsqrteLUT[12] = 16'hfe4f;
RsqrteLUT[13] = 16'hfe38;
RsqrteLUT[14] = 16'hfe23;
RsqrteLUT[15] = 16'hfe10;
RsqrteLUT[16] = 16'hfe00;
RsqrteLUT[17] = 16'hfde1;
RsqrteLUT[18] = 16'hfdc5;
RsqrteLUT[19] = 16'hfdab;
RsqrteLUT[20] = 16'hfd93;
RsqrteLUT[21] = 16'hfd7d;
RsqrteLUT[22] = 16'hfd69;
RsqrteLUT[23] = 16'hfd56;
RsqrteLUT[24] = 16'hfd44;
RsqrteLUT[25] = 16'hfd33;
RsqrteLUT[26] = 16'hfd23;
RsqrteLUT[27] = 16'hfd14;
RsqrteLUT[28] = 16'hfd06;
RsqrteLUT[29] = 16'hfcf8;
RsqrteLUT[30] = 16'hfceb;
RsqrteLUT[31] = 16'hfcdf;
RsqrteLUT[32] = 16'hfcd4;
RsqrteLUT[33] = 16'hfcc9;
RsqrteLUT[34] = 16'hfcbe;
RsqrteLUT[35] = 16'hfcb4;
RsqrteLUT[36] = 16'hfcaa;
RsqrteLUT[37] = 16'hfca1;
RsqrteLUT[38] = 16'hfc98;
RsqrteLUT[39] = 16'hfc8f;
RsqrteLUT[40] = 16'hfc87;
RsqrteLUT[41] = 16'hfc7f;
RsqrteLUT[42] = 16'hfc78;
RsqrteLUT[43] = 16'hfc70;
RsqrteLUT[44] = 16'hfc69;
RsqrteLUT[45] = 16'hfc62;
RsqrteLUT[46] = 16'hfc5b;
RsqrteLUT[47] = 16'hfc55;
RsqrteLUT[48] = 16'hfc4f;
RsqrteLUT[49] = 16'hfc49;
RsqrteLUT[50] = 16'hfc43;
RsqrteLUT[51] = 16'hfc3d;
RsqrteLUT[52] = 16'hfc38;
RsqrteLUT[53] = 16'hfc32;
RsqrteLUT[54] = 16'hfc2d;
RsqrteLUT[55] = 16'hfc28;
RsqrteLUT[56] = 16'hfc23;
RsqrteLUT[57] = 16'hfc1e;
RsqrteLUT[58] = 16'hfc19;
RsqrteLUT[59] = 16'hfc15;
RsqrteLUT[60] = 16'hfc10;
RsqrteLUT[61] = 16'hfc0c;
RsqrteLUT[62] = 16'hfc08;
RsqrteLUT[63] = 16'hfc04;
RsqrteLUT[64] = 16'hfc00;
RsqrteLUT[65] = 16'hfbf8;
RsqrteLUT[66] = 16'hfbf0;
RsqrteLUT[67] = 16'hfbe8;
RsqrteLUT[68] = 16'hfbe1;
RsqrteLUT[69] = 16'hfbda;
RsqrteLUT[70] = 16'hfbd3;
RsqrteLUT[71] = 16'hfbcc;
RsqrteLUT[72] = 16'hfbc5;
RsqrteLUT[73] = 16'hfbbe;
RsqrteLUT[74] = 16'hfbb8;
RsqrteLUT[75] = 16'hfbb1;
RsqrteLUT[76] = 16'hfbab;
RsqrteLUT[77] = 16'hfba5;
RsqrteLUT[78] = 16'hfb9f;
RsqrteLUT[79] = 16'hfb99;
RsqrteLUT[80] = 16'hfb93;
RsqrteLUT[81] = 16'hfb8e;
RsqrteLUT[82] = 16'hfb88;
RsqrteLUT[83] = 16'hfb83;
RsqrteLUT[84] = 16'hfb7d;
RsqrteLUT[85] = 16'hfb78;
RsqrteLUT[86] = 16'hfb73;
RsqrteLUT[87] = 16'hfb6e;
RsqrteLUT[88] = 16'hfb69;
RsqrteLUT[89] = 16'hfb64;
RsqrteLUT[90] = 16'hfb5f;
RsqrteLUT[91] = 16'hfb5a;
RsqrteLUT[92] = 16'hfb56;
RsqrteLUT[93] = 16'hfb51;
RsqrteLUT[94] = 16'hfb4c;
RsqrteLUT[95] = 16'hfb48;
RsqrteLUT[96] = 16'hfb44;
RsqrteLUT[97] = 16'hfb3f;
RsqrteLUT[98] = 16'hfb3b;
RsqrteLUT[99] = 16'hfb37;
RsqrteLUT[100] = 16'hfb33;
RsqrteLUT[101] = 16'hfb2f;
RsqrteLUT[102] = 16'hfb2b;
RsqrteLUT[103] = 16'hfb27;
RsqrteLUT[104] = 16'hfb23;
RsqrteLUT[105] = 16'hfb1f;
RsqrteLUT[106] = 16'hfb1b;
RsqrteLUT[107] = 16'hfb17;
RsqrteLUT[108] = 16'hfb14;
RsqrteLUT[109] = 16'hfb10;
RsqrteLUT[110] = 16'hfb0d;
RsqrteLUT[111] = 16'hfb09;
RsqrteLUT[112] = 16'hfb06;
RsqrteLUT[113] = 16'hfb02;
RsqrteLUT[114] = 16'hfaff;
RsqrteLUT[115] = 16'hfafb;
RsqrteLUT[116] = 16'hfaf8;
RsqrteLUT[117] = 16'hfaf5;
RsqrteLUT[118] = 16'hfaf2;
RsqrteLUT[119] = 16'hfaee;
RsqrteLUT[120] = 16'hfaeb;
RsqrteLUT[121] = 16'hfae8;
RsqrteLUT[122] = 16'hfae5;
RsqrteLUT[123] = 16'hfae2;
RsqrteLUT[124] = 16'hfadf;
RsqrteLUT[125] = 16'hfadc;
RsqrteLUT[126] = 16'hfad9;
RsqrteLUT[127] = 16'hfad6;
RsqrteLUT[128] = 16'hfad4;
RsqrteLUT[129] = 16'hface;
RsqrteLUT[130] = 16'hfac9;
RsqrteLUT[131] = 16'hfac3;
RsqrteLUT[132] = 16'hfabe;
RsqrteLUT[133] = 16'hfab9;
RsqrteLUT[134] = 16'hfab4;
RsqrteLUT[135] = 16'hfaaf;
RsqrteLUT[136] = 16'hfaaa;
RsqrteLUT[137] = 16'hfaa5;
RsqrteLUT[138] = 16'hfaa1;
RsqrteLUT[139] = 16'hfa9c;
RsqrteLUT[140] = 16'hfa98;
RsqrteLUT[141] = 16'hfa94;
RsqrteLUT[142] = 16'hfa8f;
RsqrteLUT[143] = 16'hfa8b;
RsqrteLUT[144] = 16'hfa87;
RsqrteLUT[145] = 16'hfa83;
RsqrteLUT[146] = 16'hfa7f;
RsqrteLUT[147] = 16'hfa7b;
RsqrteLUT[148] = 16'hfa78;
RsqrteLUT[149] = 16'hfa74;
RsqrteLUT[150] = 16'hfa70;
RsqrteLUT[151] = 16'hfa6d;
RsqrteLUT[152] = 16'hfa69;
RsqrteLUT[153] = 16'hfa66;
RsqrteLUT[154] = 16'hfa62;
RsqrteLUT[155] = 16'hfa5f;
RsqrteLUT[156] = 16'hfa5b;
RsqrteLUT[157] = 16'hfa58;
RsqrteLUT[158] = 16'hfa55;
RsqrteLUT[159] = 16'hfa52;
RsqrteLUT[160] = 16'hfa4f;
RsqrteLUT[161] = 16'hfa4c;
RsqrteLUT[162] = 16'hfa49;
RsqrteLUT[163] = 16'hfa46;
RsqrteLUT[164] = 16'hfa43;
RsqrteLUT[165] = 16'hfa40;
RsqrteLUT[166] = 16'hfa3d;
RsqrteLUT[167] = 16'hfa3a;
RsqrteLUT[168] = 16'hfa38;
RsqrteLUT[169] = 16'hfa35;
RsqrteLUT[170] = 16'hfa32;
RsqrteLUT[171] = 16'hfa2f;
RsqrteLUT[172] = 16'hfa2d;
RsqrteLUT[173] = 16'hfa2a;
RsqrteLUT[174] = 16'hfa28;
RsqrteLUT[175] = 16'hfa25;
RsqrteLUT[176] = 16'hfa23;
RsqrteLUT[177] = 16'hfa20;
RsqrteLUT[178] = 16'hfa1e;
RsqrteLUT[179] = 16'hfa1c;
RsqrteLUT[180] = 16'hfa19;
RsqrteLUT[181] = 16'hfa17;
RsqrteLUT[182] = 16'hfa15;
RsqrteLUT[183] = 16'hfa13;
RsqrteLUT[184] = 16'hfa10;
RsqrteLUT[185] = 16'hfa0e;
RsqrteLUT[186] = 16'hfa0c;
RsqrteLUT[187] = 16'hfa0a;
RsqrteLUT[188] = 16'hfa08;
RsqrteLUT[189] = 16'hfa06;
RsqrteLUT[190] = 16'hfa04;
RsqrteLUT[191] = 16'hfa02;
RsqrteLUT[192] = 16'hfa00;
RsqrteLUT[193] = 16'hf9f8;
RsqrteLUT[194] = 16'hf9f0;
RsqrteLUT[195] = 16'hf9e8;
RsqrteLUT[196] = 16'hf9e1;
RsqrteLUT[197] = 16'hf9da;
RsqrteLUT[198] = 16'hf9d3;
RsqrteLUT[199] = 16'hf9cc;
RsqrteLUT[200] = 16'hf9c5;
RsqrteLUT[201] = 16'hf9be;
RsqrteLUT[202] = 16'hf9b8;
RsqrteLUT[203] = 16'hf9b1;
RsqrteLUT[204] = 16'hf9ab;
RsqrteLUT[205] = 16'hf9a5;
RsqrteLUT[206] = 16'hf99f;
RsqrteLUT[207] = 16'hf999;
RsqrteLUT[208] = 16'hf993;
RsqrteLUT[209] = 16'hf98e;
RsqrteLUT[210] = 16'hf988;
RsqrteLUT[211] = 16'hf983;
RsqrteLUT[212] = 16'hf97d;
RsqrteLUT[213] = 16'hf978;
RsqrteLUT[214] = 16'hf973;
RsqrteLUT[215] = 16'hf96e;
RsqrteLUT[216] = 16'hf969;
RsqrteLUT[217] = 16'hf964;
RsqrteLUT[218] = 16'hf95f;
RsqrteLUT[219] = 16'hf95a;
RsqrteLUT[220] = 16'hf956;
RsqrteLUT[221] = 16'hf951;
RsqrteLUT[222] = 16'hf94c;
RsqrteLUT[223] = 16'hf948;
RsqrteLUT[224] = 16'hf944;
RsqrteLUT[225] = 16'hf93f;
RsqrteLUT[226] = 16'hf93b;
RsqrteLUT[227] = 16'hf937;
RsqrteLUT[228] = 16'hf933;
RsqrteLUT[229] = 16'hf92f;
RsqrteLUT[230] = 16'hf92b;
RsqrteLUT[231] = 16'hf927;
RsqrteLUT[232] = 16'hf923;
RsqrteLUT[233] = 16'hf91f;
RsqrteLUT[234] = 16'hf91b;
RsqrteLUT[235] = 16'hf917;
RsqrteLUT[236] = 16'hf914;
RsqrteLUT[237] = 16'hf910;
RsqrteLUT[238] = 16'hf90d;
RsqrteLUT[239] = 16'hf909;
RsqrteLUT[240] = 16'hf906;
RsqrteLUT[241] = 16'hf902;
RsqrteLUT[242] = 16'hf8ff;
RsqrteLUT[243] = 16'hf8fb;
RsqrteLUT[244] = 16'hf8f8;
RsqrteLUT[245] = 16'hf8f5;
RsqrteLUT[246] = 16'hf8f2;
RsqrteLUT[247] = 16'hf8ee;
RsqrteLUT[248] = 16'hf8eb;
RsqrteLUT[249] = 16'hf8e8;
RsqrteLUT[250] = 16'hf8e5;
RsqrteLUT[251] = 16'hf8e2;
RsqrteLUT[252] = 16'hf8df;
RsqrteLUT[253] = 16'hf8dc;
RsqrteLUT[254] = 16'hf8d9;
RsqrteLUT[255] = 16'hf8d6;
RsqrteLUT[256] = 16'hf8d4;
RsqrteLUT[257] = 16'hf8ce;
RsqrteLUT[258] = 16'hf8c9;
RsqrteLUT[259] = 16'hf8c3;
RsqrteLUT[260] = 16'hf8be;
RsqrteLUT[261] = 16'hf8b9;
RsqrteLUT[262] = 16'hf8b4;
RsqrteLUT[263] = 16'hf8af;
RsqrteLUT[264] = 16'hf8aa;
RsqrteLUT[265] = 16'hf8a5;
RsqrteLUT[266] = 16'hf8a1;
RsqrteLUT[267] = 16'hf89c;
RsqrteLUT[268] = 16'hf898;
RsqrteLUT[269] = 16'hf894;
RsqrteLUT[270] = 16'hf88f;
RsqrteLUT[271] = 16'hf88b;
RsqrteLUT[272] = 16'hf887;
RsqrteLUT[273] = 16'hf883;
RsqrteLUT[274] = 16'hf87f;
RsqrteLUT[275] = 16'hf87b;
RsqrteLUT[276] = 16'hf878;
RsqrteLUT[277] = 16'hf874;
RsqrteLUT[278] = 16'hf870;
RsqrteLUT[279] = 16'hf86d;
RsqrteLUT[280] = 16'hf869;
RsqrteLUT[281] = 16'hf866;
RsqrteLUT[282] = 16'hf862;
RsqrteLUT[283] = 16'hf85f;
RsqrteLUT[284] = 16'hf85b;
RsqrteLUT[285] = 16'hf858;
RsqrteLUT[286] = 16'hf855;
RsqrteLUT[287] = 16'hf852;
RsqrteLUT[288] = 16'hf84f;
RsqrteLUT[289] = 16'hf84c;
RsqrteLUT[290] = 16'hf849;
RsqrteLUT[291] = 16'hf846;
RsqrteLUT[292] = 16'hf843;
RsqrteLUT[293] = 16'hf840;
RsqrteLUT[294] = 16'hf83d;
RsqrteLUT[295] = 16'hf83a;
RsqrteLUT[296] = 16'hf838;
RsqrteLUT[297] = 16'hf835;
RsqrteLUT[298] = 16'hf832;
RsqrteLUT[299] = 16'hf82f;
RsqrteLUT[300] = 16'hf82d;
RsqrteLUT[301] = 16'hf82a;
RsqrteLUT[302] = 16'hf828;
RsqrteLUT[303] = 16'hf825;
RsqrteLUT[304] = 16'hf823;
RsqrteLUT[305] = 16'hf820;
RsqrteLUT[306] = 16'hf81e;
RsqrteLUT[307] = 16'hf81c;
RsqrteLUT[308] = 16'hf819;
RsqrteLUT[309] = 16'hf817;
RsqrteLUT[310] = 16'hf815;
RsqrteLUT[311] = 16'hf813;
RsqrteLUT[312] = 16'hf810;
RsqrteLUT[313] = 16'hf80e;
RsqrteLUT[314] = 16'hf80c;
RsqrteLUT[315] = 16'hf80a;
RsqrteLUT[316] = 16'hf808;
RsqrteLUT[317] = 16'hf806;
RsqrteLUT[318] = 16'hf804;
RsqrteLUT[319] = 16'hf802;
RsqrteLUT[320] = 16'hf800;
RsqrteLUT[321] = 16'hf7f8;
RsqrteLUT[322] = 16'hf7f0;
RsqrteLUT[323] = 16'hf7e8;
RsqrteLUT[324] = 16'hf7e1;
RsqrteLUT[325] = 16'hf7da;
RsqrteLUT[326] = 16'hf7d3;
RsqrteLUT[327] = 16'hf7cc;
RsqrteLUT[328] = 16'hf7c5;
RsqrteLUT[329] = 16'hf7be;
RsqrteLUT[330] = 16'hf7b8;
RsqrteLUT[331] = 16'hf7b1;
RsqrteLUT[332] = 16'hf7ab;
RsqrteLUT[333] = 16'hf7a5;
RsqrteLUT[334] = 16'hf79f;
RsqrteLUT[335] = 16'hf799;
RsqrteLUT[336] = 16'hf793;
RsqrteLUT[337] = 16'hf78e;
RsqrteLUT[338] = 16'hf788;
RsqrteLUT[339] = 16'hf783;
RsqrteLUT[340] = 16'hf77d;
RsqrteLUT[341] = 16'hf778;
RsqrteLUT[342] = 16'hf773;
RsqrteLUT[343] = 16'hf76e;
RsqrteLUT[344] = 16'hf769;
RsqrteLUT[345] = 16'hf764;
RsqrteLUT[346] = 16'hf75f;
RsqrteLUT[347] = 16'hf75a;
RsqrteLUT[348] = 16'hf756;
RsqrteLUT[349] = 16'hf751;
RsqrteLUT[350] = 16'hf74c;
RsqrteLUT[351] = 16'hf748;
RsqrteLUT[352] = 16'hf744;
RsqrteLUT[353] = 16'hf73f;
RsqrteLUT[354] = 16'hf73b;
RsqrteLUT[355] = 16'hf737;
RsqrteLUT[356] = 16'hf733;
RsqrteLUT[357] = 16'hf72f;
RsqrteLUT[358] = 16'hf72b;
RsqrteLUT[359] = 16'hf727;
RsqrteLUT[360] = 16'hf723;
RsqrteLUT[361] = 16'hf71f;
RsqrteLUT[362] = 16'hf71b;
RsqrteLUT[363] = 16'hf717;
RsqrteLUT[364] = 16'hf714;
RsqrteLUT[365] = 16'hf710;
RsqrteLUT[366] = 16'hf70d;
RsqrteLUT[367] = 16'hf709;
RsqrteLUT[368] = 16'hf706;
RsqrteLUT[369] = 16'hf702;
RsqrteLUT[370] = 16'hf6ff;
RsqrteLUT[371] = 16'hf6fb;
RsqrteLUT[372] = 16'hf6f8;
RsqrteLUT[373] = 16'hf6f5;
RsqrteLUT[374] = 16'hf6f2;
RsqrteLUT[375] = 16'hf6ee;
RsqrteLUT[376] = 16'hf6eb;
RsqrteLUT[377] = 16'hf6e8;
RsqrteLUT[378] = 16'hf6e5;
RsqrteLUT[379] = 16'hf6e2;
RsqrteLUT[380] = 16'hf6df;
RsqrteLUT[381] = 16'hf6dc;
RsqrteLUT[382] = 16'hf6d9;
RsqrteLUT[383] = 16'hf6d6;
RsqrteLUT[384] = 16'hf6d4;
RsqrteLUT[385] = 16'hf6ce;
RsqrteLUT[386] = 16'hf6c9;
RsqrteLUT[387] = 16'hf6c3;
RsqrteLUT[388] = 16'hf6be;
RsqrteLUT[389] = 16'hf6b9;
RsqrteLUT[390] = 16'hf6b4;
RsqrteLUT[391] = 16'hf6af;
RsqrteLUT[392] = 16'hf6aa;
RsqrteLUT[393] = 16'hf6a5;
RsqrteLUT[394] = 16'hf6a1;
RsqrteLUT[395] = 16'hf69c;
RsqrteLUT[396] = 16'hf698;
RsqrteLUT[397] = 16'hf694;
RsqrteLUT[398] = 16'hf68f;
RsqrteLUT[399] = 16'hf68b;
RsqrteLUT[400] = 16'hf687;
RsqrteLUT[401] = 16'hf683;
RsqrteLUT[402] = 16'hf67f;
RsqrteLUT[403] = 16'hf67b;
RsqrteLUT[404] = 16'hf678;
RsqrteLUT[405] = 16'hf674;
RsqrteLUT[406] = 16'hf670;
RsqrteLUT[407] = 16'hf66d;
RsqrteLUT[408] = 16'hf669;
RsqrteLUT[409] = 16'hf666;
RsqrteLUT[410] = 16'hf662;
RsqrteLUT[411] = 16'hf65f;
RsqrteLUT[412] = 16'hf65b;
RsqrteLUT[413] = 16'hf658;
RsqrteLUT[414] = 16'hf655;
RsqrteLUT[415] = 16'hf652;
RsqrteLUT[416] = 16'hf64f;
RsqrteLUT[417] = 16'hf64c;
RsqrteLUT[418] = 16'hf649;
RsqrteLUT[419] = 16'hf646;
RsqrteLUT[420] = 16'hf643;
RsqrteLUT[421] = 16'hf640;
RsqrteLUT[422] = 16'hf63d;
RsqrteLUT[423] = 16'hf63a;
RsqrteLUT[424] = 16'hf638;
RsqrteLUT[425] = 16'hf635;
RsqrteLUT[426] = 16'hf632;
RsqrteLUT[427] = 16'hf62f;
RsqrteLUT[428] = 16'hf62d;
RsqrteLUT[429] = 16'hf62a;
RsqrteLUT[430] = 16'hf628;
RsqrteLUT[431] = 16'hf625;
RsqrteLUT[432] = 16'hf623;
RsqrteLUT[433] = 16'hf620;
RsqrteLUT[434] = 16'hf61e;
RsqrteLUT[435] = 16'hf61c;
RsqrteLUT[436] = 16'hf619;
RsqrteLUT[437] = 16'hf617;
RsqrteLUT[438] = 16'hf615;
RsqrteLUT[439] = 16'hf613;
RsqrteLUT[440] = 16'hf610;
RsqrteLUT[441] = 16'hf60e;
RsqrteLUT[442] = 16'hf60c;
RsqrteLUT[443] = 16'hf60a;
RsqrteLUT[444] = 16'hf608;
RsqrteLUT[445] = 16'hf606;
RsqrteLUT[446] = 16'hf604;
RsqrteLUT[447] = 16'hf602;
RsqrteLUT[448] = 16'hf600;
RsqrteLUT[449] = 16'hf5f8;
RsqrteLUT[450] = 16'hf5f0;
RsqrteLUT[451] = 16'hf5e8;
RsqrteLUT[452] = 16'hf5e1;
RsqrteLUT[453] = 16'hf5da;
RsqrteLUT[454] = 16'hf5d3;
RsqrteLUT[455] = 16'hf5cc;
RsqrteLUT[456] = 16'hf5c5;
RsqrteLUT[457] = 16'hf5be;
RsqrteLUT[458] = 16'hf5b8;
RsqrteLUT[459] = 16'hf5b1;
RsqrteLUT[460] = 16'hf5ab;
RsqrteLUT[461] = 16'hf5a5;
RsqrteLUT[462] = 16'hf59f;
RsqrteLUT[463] = 16'hf599;
RsqrteLUT[464] = 16'hf593;
RsqrteLUT[465] = 16'hf58e;
RsqrteLUT[466] = 16'hf588;
RsqrteLUT[467] = 16'hf583;
RsqrteLUT[468] = 16'hf57d;
RsqrteLUT[469] = 16'hf578;
RsqrteLUT[470] = 16'hf573;
RsqrteLUT[471] = 16'hf56e;
RsqrteLUT[472] = 16'hf569;
RsqrteLUT[473] = 16'hf564;
RsqrteLUT[474] = 16'hf55f;
RsqrteLUT[475] = 16'hf55a;
RsqrteLUT[476] = 16'hf556;
RsqrteLUT[477] = 16'hf551;
RsqrteLUT[478] = 16'hf54c;
RsqrteLUT[479] = 16'hf548;
RsqrteLUT[480] = 16'hf544;
RsqrteLUT[481] = 16'hf53f;
RsqrteLUT[482] = 16'hf53b;
RsqrteLUT[483] = 16'hf537;
RsqrteLUT[484] = 16'hf533;
RsqrteLUT[485] = 16'hf52f;
RsqrteLUT[486] = 16'hf52b;
RsqrteLUT[487] = 16'hf527;
RsqrteLUT[488] = 16'hf523;
RsqrteLUT[489] = 16'hf51f;
RsqrteLUT[490] = 16'hf51b;
RsqrteLUT[491] = 16'hf517;
RsqrteLUT[492] = 16'hf514;
RsqrteLUT[493] = 16'hf510;
RsqrteLUT[494] = 16'hf50d;
RsqrteLUT[495] = 16'hf509;
RsqrteLUT[496] = 16'hf506;
RsqrteLUT[497] = 16'hf502;
RsqrteLUT[498] = 16'hf4ff;
RsqrteLUT[499] = 16'hf4fb;
RsqrteLUT[500] = 16'hf4f8;
RsqrteLUT[501] = 16'hf4f5;
RsqrteLUT[502] = 16'hf4f2;
RsqrteLUT[503] = 16'hf4ee;
RsqrteLUT[504] = 16'hf4eb;
RsqrteLUT[505] = 16'hf4e8;
RsqrteLUT[506] = 16'hf4e5;
RsqrteLUT[507] = 16'hf4e2;
RsqrteLUT[508] = 16'hf4df;
RsqrteLUT[509] = 16'hf4dc;
RsqrteLUT[510] = 16'hf4d9;
RsqrteLUT[511] = 16'hf4d6;
RsqrteLUT[512] = 16'hf4d4;
RsqrteLUT[513] = 16'hf4ce;
RsqrteLUT[514] = 16'hf4c9;
RsqrteLUT[515] = 16'hf4c3;
RsqrteLUT[516] = 16'hf4be;
RsqrteLUT[517] = 16'hf4b9;
RsqrteLUT[518] = 16'hf4b4;
RsqrteLUT[519] = 16'hf4af;
RsqrteLUT[520] = 16'hf4aa;
RsqrteLUT[521] = 16'hf4a5;
RsqrteLUT[522] = 16'hf4a1;
RsqrteLUT[523] = 16'hf49c;
RsqrteLUT[524] = 16'hf498;
RsqrteLUT[525] = 16'hf494;
RsqrteLUT[526] = 16'hf48f;
RsqrteLUT[527] = 16'hf48b;
RsqrteLUT[528] = 16'hf487;
RsqrteLUT[529] = 16'hf483;
RsqrteLUT[530] = 16'hf47f;
RsqrteLUT[531] = 16'hf47b;
RsqrteLUT[532] = 16'hf478;
RsqrteLUT[533] = 16'hf474;
RsqrteLUT[534] = 16'hf470;
RsqrteLUT[535] = 16'hf46d;
RsqrteLUT[536] = 16'hf469;
RsqrteLUT[537] = 16'hf466;
RsqrteLUT[538] = 16'hf462;
RsqrteLUT[539] = 16'hf45f;
RsqrteLUT[540] = 16'hf45b;
RsqrteLUT[541] = 16'hf458;
RsqrteLUT[542] = 16'hf455;
RsqrteLUT[543] = 16'hf452;
RsqrteLUT[544] = 16'hf44f;
RsqrteLUT[545] = 16'hf44c;
RsqrteLUT[546] = 16'hf449;
RsqrteLUT[547] = 16'hf446;
RsqrteLUT[548] = 16'hf443;
RsqrteLUT[549] = 16'hf440;
RsqrteLUT[550] = 16'hf43d;
RsqrteLUT[551] = 16'hf43a;
RsqrteLUT[552] = 16'hf438;
RsqrteLUT[553] = 16'hf435;
RsqrteLUT[554] = 16'hf432;
RsqrteLUT[555] = 16'hf42f;
RsqrteLUT[556] = 16'hf42d;
RsqrteLUT[557] = 16'hf42a;
RsqrteLUT[558] = 16'hf428;
RsqrteLUT[559] = 16'hf425;
RsqrteLUT[560] = 16'hf423;
RsqrteLUT[561] = 16'hf420;
RsqrteLUT[562] = 16'hf41e;
RsqrteLUT[563] = 16'hf41c;
RsqrteLUT[564] = 16'hf419;
RsqrteLUT[565] = 16'hf417;
RsqrteLUT[566] = 16'hf415;
RsqrteLUT[567] = 16'hf413;
RsqrteLUT[568] = 16'hf410;
RsqrteLUT[569] = 16'hf40e;
RsqrteLUT[570] = 16'hf40c;
RsqrteLUT[571] = 16'hf40a;
RsqrteLUT[572] = 16'hf408;
RsqrteLUT[573] = 16'hf406;
RsqrteLUT[574] = 16'hf404;
RsqrteLUT[575] = 16'hf402;
RsqrteLUT[576] = 16'hf400;
RsqrteLUT[577] = 16'hf3f8;
RsqrteLUT[578] = 16'hf3f0;
RsqrteLUT[579] = 16'hf3e8;
RsqrteLUT[580] = 16'hf3e1;
RsqrteLUT[581] = 16'hf3da;
RsqrteLUT[582] = 16'hf3d3;
RsqrteLUT[583] = 16'hf3cc;
RsqrteLUT[584] = 16'hf3c5;
RsqrteLUT[585] = 16'hf3be;
RsqrteLUT[586] = 16'hf3b8;
RsqrteLUT[587] = 16'hf3b1;
RsqrteLUT[588] = 16'hf3ab;
RsqrteLUT[589] = 16'hf3a5;
RsqrteLUT[590] = 16'hf39f;
RsqrteLUT[591] = 16'hf399;
RsqrteLUT[592] = 16'hf393;
RsqrteLUT[593] = 16'hf38e;
RsqrteLUT[594] = 16'hf388;
RsqrteLUT[595] = 16'hf383;
RsqrteLUT[596] = 16'hf37d;
RsqrteLUT[597] = 16'hf378;
RsqrteLUT[598] = 16'hf373;
RsqrteLUT[599] = 16'hf36e;
RsqrteLUT[600] = 16'hf369;
RsqrteLUT[601] = 16'hf364;
RsqrteLUT[602] = 16'hf35f;
RsqrteLUT[603] = 16'hf35a;
RsqrteLUT[604] = 16'hf356;
RsqrteLUT[605] = 16'hf351;
RsqrteLUT[606] = 16'hf34c;
RsqrteLUT[607] = 16'hf348;
RsqrteLUT[608] = 16'hf344;
RsqrteLUT[609] = 16'hf33f;
RsqrteLUT[610] = 16'hf33b;
RsqrteLUT[611] = 16'hf337;
RsqrteLUT[612] = 16'hf333;
RsqrteLUT[613] = 16'hf32f;
RsqrteLUT[614] = 16'hf32b;
RsqrteLUT[615] = 16'hf327;
RsqrteLUT[616] = 16'hf323;
RsqrteLUT[617] = 16'hf31f;
RsqrteLUT[618] = 16'hf31b;
RsqrteLUT[619] = 16'hf317;
RsqrteLUT[620] = 16'hf314;
RsqrteLUT[621] = 16'hf310;
RsqrteLUT[622] = 16'hf30d;
RsqrteLUT[623] = 16'hf309;
RsqrteLUT[624] = 16'hf306;
RsqrteLUT[625] = 16'hf302;
RsqrteLUT[626] = 16'hf2ff;
RsqrteLUT[627] = 16'hf2fb;
RsqrteLUT[628] = 16'hf2f8;
RsqrteLUT[629] = 16'hf2f5;
RsqrteLUT[630] = 16'hf2f2;
RsqrteLUT[631] = 16'hf2ee;
RsqrteLUT[632] = 16'hf2eb;
RsqrteLUT[633] = 16'hf2e8;
RsqrteLUT[634] = 16'hf2e5;
RsqrteLUT[635] = 16'hf2e2;
RsqrteLUT[636] = 16'hf2df;
RsqrteLUT[637] = 16'hf2dc;
RsqrteLUT[638] = 16'hf2d9;
RsqrteLUT[639] = 16'hf2d6;
RsqrteLUT[640] = 16'hf2d4;
RsqrteLUT[641] = 16'hf2ce;
RsqrteLUT[642] = 16'hf2c9;
RsqrteLUT[643] = 16'hf2c3;
RsqrteLUT[644] = 16'hf2be;
RsqrteLUT[645] = 16'hf2b9;
RsqrteLUT[646] = 16'hf2b4;
RsqrteLUT[647] = 16'hf2af;
RsqrteLUT[648] = 16'hf2aa;
RsqrteLUT[649] = 16'hf2a5;
RsqrteLUT[650] = 16'hf2a1;
RsqrteLUT[651] = 16'hf29c;
RsqrteLUT[652] = 16'hf298;
RsqrteLUT[653] = 16'hf294;
RsqrteLUT[654] = 16'hf28f;
RsqrteLUT[655] = 16'hf28b;
RsqrteLUT[656] = 16'hf287;
RsqrteLUT[657] = 16'hf283;
RsqrteLUT[658] = 16'hf27f;
RsqrteLUT[659] = 16'hf27b;
RsqrteLUT[660] = 16'hf278;
RsqrteLUT[661] = 16'hf274;
RsqrteLUT[662] = 16'hf270;
RsqrteLUT[663] = 16'hf26d;
RsqrteLUT[664] = 16'hf269;
RsqrteLUT[665] = 16'hf266;
RsqrteLUT[666] = 16'hf262;
RsqrteLUT[667] = 16'hf25f;
RsqrteLUT[668] = 16'hf25b;
RsqrteLUT[669] = 16'hf258;
RsqrteLUT[670] = 16'hf255;
RsqrteLUT[671] = 16'hf252;
RsqrteLUT[672] = 16'hf24f;
RsqrteLUT[673] = 16'hf24c;
RsqrteLUT[674] = 16'hf249;
RsqrteLUT[675] = 16'hf246;
RsqrteLUT[676] = 16'hf243;
RsqrteLUT[677] = 16'hf240;
RsqrteLUT[678] = 16'hf23d;
RsqrteLUT[679] = 16'hf23a;
RsqrteLUT[680] = 16'hf238;
RsqrteLUT[681] = 16'hf235;
RsqrteLUT[682] = 16'hf232;
RsqrteLUT[683] = 16'hf22f;
RsqrteLUT[684] = 16'hf22d;
RsqrteLUT[685] = 16'hf22a;
RsqrteLUT[686] = 16'hf228;
RsqrteLUT[687] = 16'hf225;
RsqrteLUT[688] = 16'hf223;
RsqrteLUT[689] = 16'hf220;
RsqrteLUT[690] = 16'hf21e;
RsqrteLUT[691] = 16'hf21c;
RsqrteLUT[692] = 16'hf219;
RsqrteLUT[693] = 16'hf217;
RsqrteLUT[694] = 16'hf215;
RsqrteLUT[695] = 16'hf213;
RsqrteLUT[696] = 16'hf210;
RsqrteLUT[697] = 16'hf20e;
RsqrteLUT[698] = 16'hf20c;
RsqrteLUT[699] = 16'hf20a;
RsqrteLUT[700] = 16'hf208;
RsqrteLUT[701] = 16'hf206;
RsqrteLUT[702] = 16'hf204;
RsqrteLUT[703] = 16'hf202;
RsqrteLUT[704] = 16'hf200;
RsqrteLUT[705] = 16'hf1f8;
RsqrteLUT[706] = 16'hf1f0;
RsqrteLUT[707] = 16'hf1e8;
RsqrteLUT[708] = 16'hf1e1;
RsqrteLUT[709] = 16'hf1da;
RsqrteLUT[710] = 16'hf1d3;
RsqrteLUT[711] = 16'hf1cc;
RsqrteLUT[712] = 16'hf1c5;
RsqrteLUT[713] = 16'hf1be;
RsqrteLUT[714] = 16'hf1b8;
RsqrteLUT[715] = 16'hf1b1;
RsqrteLUT[716] = 16'hf1ab;
RsqrteLUT[717] = 16'hf1a5;
RsqrteLUT[718] = 16'hf19f;
RsqrteLUT[719] = 16'hf199;
RsqrteLUT[720] = 16'hf193;
RsqrteLUT[721] = 16'hf18e;
RsqrteLUT[722] = 16'hf188;
RsqrteLUT[723] = 16'hf183;
RsqrteLUT[724] = 16'hf17d;
RsqrteLUT[725] = 16'hf178;
RsqrteLUT[726] = 16'hf173;
RsqrteLUT[727] = 16'hf16e;
RsqrteLUT[728] = 16'hf169;
RsqrteLUT[729] = 16'hf164;
RsqrteLUT[730] = 16'hf15f;
RsqrteLUT[731] = 16'hf15a;
RsqrteLUT[732] = 16'hf156;
RsqrteLUT[733] = 16'hf151;
RsqrteLUT[734] = 16'hf14c;
RsqrteLUT[735] = 16'hf148;
RsqrteLUT[736] = 16'hf144;
RsqrteLUT[737] = 16'hf13f;
RsqrteLUT[738] = 16'hf13b;
RsqrteLUT[739] = 16'hf137;
RsqrteLUT[740] = 16'hf133;
RsqrteLUT[741] = 16'hf12f;
RsqrteLUT[742] = 16'hf12b;
RsqrteLUT[743] = 16'hf127;
RsqrteLUT[744] = 16'hf123;
RsqrteLUT[745] = 16'hf11f;
RsqrteLUT[746] = 16'hf11b;
RsqrteLUT[747] = 16'hf117;
RsqrteLUT[748] = 16'hf114;
RsqrteLUT[749] = 16'hf110;
RsqrteLUT[750] = 16'hf10d;
RsqrteLUT[751] = 16'hf109;
RsqrteLUT[752] = 16'hf106;
RsqrteLUT[753] = 16'hf102;
RsqrteLUT[754] = 16'hf0ff;
RsqrteLUT[755] = 16'hf0fb;
RsqrteLUT[756] = 16'hf0f8;
RsqrteLUT[757] = 16'hf0f5;
RsqrteLUT[758] = 16'hf0f2;
RsqrteLUT[759] = 16'hf0ee;
RsqrteLUT[760] = 16'hf0eb;
RsqrteLUT[761] = 16'hf0e8;
RsqrteLUT[762] = 16'hf0e5;
RsqrteLUT[763] = 16'hf0e2;
RsqrteLUT[764] = 16'hf0df;
RsqrteLUT[765] = 16'hf0dc;
RsqrteLUT[766] = 16'hf0d9;
RsqrteLUT[767] = 16'hf0d6;
RsqrteLUT[768] = 16'hf0d4;
RsqrteLUT[769] = 16'hf0ce;
RsqrteLUT[770] = 16'hf0c9;
RsqrteLUT[771] = 16'hf0c3;
RsqrteLUT[772] = 16'hf0be;
RsqrteLUT[773] = 16'hf0b9;
RsqrteLUT[774] = 16'hf0b4;
RsqrteLUT[775] = 16'hf0af;
RsqrteLUT[776] = 16'hf0aa;
RsqrteLUT[777] = 16'hf0a5;
RsqrteLUT[778] = 16'hf0a1;
RsqrteLUT[779] = 16'hf09c;
RsqrteLUT[780] = 16'hf098;
RsqrteLUT[781] = 16'hf094;
RsqrteLUT[782] = 16'hf08f;
RsqrteLUT[783] = 16'hf08b;
RsqrteLUT[784] = 16'hf087;
RsqrteLUT[785] = 16'hf083;
RsqrteLUT[786] = 16'hf07f;
RsqrteLUT[787] = 16'hf07b;
RsqrteLUT[788] = 16'hf078;
RsqrteLUT[789] = 16'hf074;
RsqrteLUT[790] = 16'hf070;
RsqrteLUT[791] = 16'hf06d;
RsqrteLUT[792] = 16'hf069;
RsqrteLUT[793] = 16'hf066;
RsqrteLUT[794] = 16'hf062;
RsqrteLUT[795] = 16'hf05f;
RsqrteLUT[796] = 16'hf05b;
RsqrteLUT[797] = 16'hf058;
RsqrteLUT[798] = 16'hf055;
RsqrteLUT[799] = 16'hf052;
RsqrteLUT[800] = 16'hf04f;
RsqrteLUT[801] = 16'hf04c;
RsqrteLUT[802] = 16'hf049;
RsqrteLUT[803] = 16'hf046;
RsqrteLUT[804] = 16'hf043;
RsqrteLUT[805] = 16'hf040;
RsqrteLUT[806] = 16'hf03d;
RsqrteLUT[807] = 16'hf03a;
RsqrteLUT[808] = 16'hf038;
RsqrteLUT[809] = 16'hf035;
RsqrteLUT[810] = 16'hf032;
RsqrteLUT[811] = 16'hf02f;
RsqrteLUT[812] = 16'hf02d;
RsqrteLUT[813] = 16'hf02a;
RsqrteLUT[814] = 16'hf028;
RsqrteLUT[815] = 16'hf025;
RsqrteLUT[816] = 16'hf023;
RsqrteLUT[817] = 16'hf020;
RsqrteLUT[818] = 16'hf01e;
RsqrteLUT[819] = 16'hf01c;
RsqrteLUT[820] = 16'hf019;
RsqrteLUT[821] = 16'hf017;
RsqrteLUT[822] = 16'hf015;
RsqrteLUT[823] = 16'hf013;
RsqrteLUT[824] = 16'hf010;
RsqrteLUT[825] = 16'hf00e;
RsqrteLUT[826] = 16'hf00c;
RsqrteLUT[827] = 16'hf00a;
RsqrteLUT[828] = 16'hf008;
RsqrteLUT[829] = 16'hf006;
RsqrteLUT[830] = 16'hf004;
RsqrteLUT[831] = 16'hf002;
RsqrteLUT[832] = 16'hf000;
RsqrteLUT[833] = 16'heff8;
RsqrteLUT[834] = 16'heff0;
RsqrteLUT[835] = 16'hefe8;
RsqrteLUT[836] = 16'hefe1;
RsqrteLUT[837] = 16'hefda;
RsqrteLUT[838] = 16'hefd3;
RsqrteLUT[839] = 16'hefcc;
RsqrteLUT[840] = 16'hefc5;
RsqrteLUT[841] = 16'hefbe;
RsqrteLUT[842] = 16'hefb8;
RsqrteLUT[843] = 16'hefb1;
RsqrteLUT[844] = 16'hefab;
RsqrteLUT[845] = 16'hefa5;
RsqrteLUT[846] = 16'hef9f;
RsqrteLUT[847] = 16'hef99;
RsqrteLUT[848] = 16'hef93;
RsqrteLUT[849] = 16'hef8e;
RsqrteLUT[850] = 16'hef88;
RsqrteLUT[851] = 16'hef83;
RsqrteLUT[852] = 16'hef7d;
RsqrteLUT[853] = 16'hef78;
RsqrteLUT[854] = 16'hef73;
RsqrteLUT[855] = 16'hef6e;
RsqrteLUT[856] = 16'hef69;
RsqrteLUT[857] = 16'hef64;
RsqrteLUT[858] = 16'hef5f;
RsqrteLUT[859] = 16'hef5a;
RsqrteLUT[860] = 16'hef56;
RsqrteLUT[861] = 16'hef51;
RsqrteLUT[862] = 16'hef4c;
RsqrteLUT[863] = 16'hef48;
RsqrteLUT[864] = 16'hef44;
RsqrteLUT[865] = 16'hef3f;
RsqrteLUT[866] = 16'hef3b;
RsqrteLUT[867] = 16'hef37;
RsqrteLUT[868] = 16'hef33;
RsqrteLUT[869] = 16'hef2f;
RsqrteLUT[870] = 16'hef2b;
RsqrteLUT[871] = 16'hef27;
RsqrteLUT[872] = 16'hef23;
RsqrteLUT[873] = 16'hef1f;
RsqrteLUT[874] = 16'hef1b;
RsqrteLUT[875] = 16'hef17;
RsqrteLUT[876] = 16'hef14;
RsqrteLUT[877] = 16'hef10;
RsqrteLUT[878] = 16'hef0d;
RsqrteLUT[879] = 16'hef09;
RsqrteLUT[880] = 16'hef06;
RsqrteLUT[881] = 16'hef02;
RsqrteLUT[882] = 16'heeff;
RsqrteLUT[883] = 16'heefb;
RsqrteLUT[884] = 16'heef8;
RsqrteLUT[885] = 16'heef5;
RsqrteLUT[886] = 16'heef2;
RsqrteLUT[887] = 16'heeee;
RsqrteLUT[888] = 16'heeeb;
RsqrteLUT[889] = 16'heee8;
RsqrteLUT[890] = 16'heee5;
RsqrteLUT[891] = 16'heee2;
RsqrteLUT[892] = 16'heedf;
RsqrteLUT[893] = 16'heedc;
RsqrteLUT[894] = 16'heed9;
RsqrteLUT[895] = 16'heed6;
RsqrteLUT[896] = 16'heed4;
RsqrteLUT[897] = 16'heece;
RsqrteLUT[898] = 16'heec9;
RsqrteLUT[899] = 16'heec3;
RsqrteLUT[900] = 16'heebe;
RsqrteLUT[901] = 16'heeb9;
RsqrteLUT[902] = 16'heeb4;
RsqrteLUT[903] = 16'heeaf;
RsqrteLUT[904] = 16'heeaa;
RsqrteLUT[905] = 16'heea5;
RsqrteLUT[906] = 16'heea1;
RsqrteLUT[907] = 16'hee9c;
RsqrteLUT[908] = 16'hee98;
RsqrteLUT[909] = 16'hee94;
RsqrteLUT[910] = 16'hee8f;
RsqrteLUT[911] = 16'hee8b;
RsqrteLUT[912] = 16'hee87;
RsqrteLUT[913] = 16'hee83;
RsqrteLUT[914] = 16'hee7f;
RsqrteLUT[915] = 16'hee7b;
RsqrteLUT[916] = 16'hee78;
RsqrteLUT[917] = 16'hee74;
RsqrteLUT[918] = 16'hee70;
RsqrteLUT[919] = 16'hee6d;
RsqrteLUT[920] = 16'hee69;
RsqrteLUT[921] = 16'hee66;
RsqrteLUT[922] = 16'hee62;
RsqrteLUT[923] = 16'hee5f;
RsqrteLUT[924] = 16'hee5b;
RsqrteLUT[925] = 16'hee58;
RsqrteLUT[926] = 16'hee55;
RsqrteLUT[927] = 16'hee52;
RsqrteLUT[928] = 16'hee4f;
RsqrteLUT[929] = 16'hee4c;
RsqrteLUT[930] = 16'hee49;
RsqrteLUT[931] = 16'hee46;
RsqrteLUT[932] = 16'hee43;
RsqrteLUT[933] = 16'hee40;
RsqrteLUT[934] = 16'hee3d;
RsqrteLUT[935] = 16'hee3a;
RsqrteLUT[936] = 16'hee38;
RsqrteLUT[937] = 16'hee35;
RsqrteLUT[938] = 16'hee32;
RsqrteLUT[939] = 16'hee2f;
RsqrteLUT[940] = 16'hee2d;
RsqrteLUT[941] = 16'hee2a;
RsqrteLUT[942] = 16'hee28;
RsqrteLUT[943] = 16'hee25;
RsqrteLUT[944] = 16'hee23;
RsqrteLUT[945] = 16'hee20;
RsqrteLUT[946] = 16'hee1e;
RsqrteLUT[947] = 16'hee1c;
RsqrteLUT[948] = 16'hee19;
RsqrteLUT[949] = 16'hee17;
RsqrteLUT[950] = 16'hee15;
RsqrteLUT[951] = 16'hee13;
RsqrteLUT[952] = 16'hee10;
RsqrteLUT[953] = 16'hee0e;
RsqrteLUT[954] = 16'hee0c;
RsqrteLUT[955] = 16'hee0a;
RsqrteLUT[956] = 16'hee08;
RsqrteLUT[957] = 16'hee06;
RsqrteLUT[958] = 16'hee04;
RsqrteLUT[959] = 16'hee02;
RsqrteLUT[960] = 16'hee00;
RsqrteLUT[961] = 16'hedf8;
RsqrteLUT[962] = 16'hedf0;
RsqrteLUT[963] = 16'hede8;
RsqrteLUT[964] = 16'hede1;
RsqrteLUT[965] = 16'hedda;
RsqrteLUT[966] = 16'hedd3;
RsqrteLUT[967] = 16'hedcc;
RsqrteLUT[968] = 16'hedc5;
RsqrteLUT[969] = 16'hedbe;
RsqrteLUT[970] = 16'hedb8;
RsqrteLUT[971] = 16'hedb1;
RsqrteLUT[972] = 16'hedab;
RsqrteLUT[973] = 16'heda5;
RsqrteLUT[974] = 16'hed9f;
RsqrteLUT[975] = 16'hed99;
RsqrteLUT[976] = 16'hed93;
RsqrteLUT[977] = 16'hed8e;
RsqrteLUT[978] = 16'hed88;
RsqrteLUT[979] = 16'hed83;
RsqrteLUT[980] = 16'hed7d;
RsqrteLUT[981] = 16'hed78;
RsqrteLUT[982] = 16'hed73;
RsqrteLUT[983] = 16'hed6e;
RsqrteLUT[984] = 16'hed69;
RsqrteLUT[985] = 16'hed64;
RsqrteLUT[986] = 16'hed5f;
RsqrteLUT[987] = 16'hed5a;
RsqrteLUT[988] = 16'hed56;
RsqrteLUT[989] = 16'hed51;
RsqrteLUT[990] = 16'hed4c;
RsqrteLUT[991] = 16'hed48;
RsqrteLUT[992] = 16'hed44;
RsqrteLUT[993] = 16'hed3f;
RsqrteLUT[994] = 16'hed3b;
RsqrteLUT[995] = 16'hed37;
RsqrteLUT[996] = 16'hed33;
RsqrteLUT[997] = 16'hed2f;
RsqrteLUT[998] = 16'hed2b;
RsqrteLUT[999] = 16'hed27;
RsqrteLUT[1000] = 16'hed23;
RsqrteLUT[1001] = 16'hed1f;
RsqrteLUT[1002] = 16'hed1b;
RsqrteLUT[1003] = 16'hed17;
RsqrteLUT[1004] = 16'hed14;
RsqrteLUT[1005] = 16'hed10;
RsqrteLUT[1006] = 16'hed0d;
RsqrteLUT[1007] = 16'hed09;
RsqrteLUT[1008] = 16'hed06;
RsqrteLUT[1009] = 16'hed02;
RsqrteLUT[1010] = 16'hecff;
RsqrteLUT[1011] = 16'hecfb;
RsqrteLUT[1012] = 16'hecf8;
RsqrteLUT[1013] = 16'hecf5;
RsqrteLUT[1014] = 16'hecf2;
RsqrteLUT[1015] = 16'hecee;
RsqrteLUT[1016] = 16'heceb;
RsqrteLUT[1017] = 16'hece8;
RsqrteLUT[1018] = 16'hece5;
RsqrteLUT[1019] = 16'hece2;
RsqrteLUT[1020] = 16'hecdf;
RsqrteLUT[1021] = 16'hecdc;
RsqrteLUT[1022] = 16'hecd9;
RsqrteLUT[1023] = 16'hecd6;
RsqrteLUT[1024] = 16'hecd4;
RsqrteLUT[1025] = 16'hecce;
RsqrteLUT[1026] = 16'hecc9;
RsqrteLUT[1027] = 16'hecc3;
RsqrteLUT[1028] = 16'hecbe;
RsqrteLUT[1029] = 16'hecb9;
RsqrteLUT[1030] = 16'hecb4;
RsqrteLUT[1031] = 16'hecaf;
RsqrteLUT[1032] = 16'hecaa;
RsqrteLUT[1033] = 16'heca5;
RsqrteLUT[1034] = 16'heca1;
RsqrteLUT[1035] = 16'hec9c;
RsqrteLUT[1036] = 16'hec98;
RsqrteLUT[1037] = 16'hec94;
RsqrteLUT[1038] = 16'hec8f;
RsqrteLUT[1039] = 16'hec8b;
RsqrteLUT[1040] = 16'hec87;
RsqrteLUT[1041] = 16'hec83;
RsqrteLUT[1042] = 16'hec7f;
RsqrteLUT[1043] = 16'hec7b;
RsqrteLUT[1044] = 16'hec78;
RsqrteLUT[1045] = 16'hec74;
RsqrteLUT[1046] = 16'hec70;
RsqrteLUT[1047] = 16'hec6d;
RsqrteLUT[1048] = 16'hec69;
RsqrteLUT[1049] = 16'hec66;
RsqrteLUT[1050] = 16'hec62;
RsqrteLUT[1051] = 16'hec5f;
RsqrteLUT[1052] = 16'hec5b;
RsqrteLUT[1053] = 16'hec58;
RsqrteLUT[1054] = 16'hec55;
RsqrteLUT[1055] = 16'hec52;
RsqrteLUT[1056] = 16'hec4f;
RsqrteLUT[1057] = 16'hec4c;
RsqrteLUT[1058] = 16'hec49;
RsqrteLUT[1059] = 16'hec46;
RsqrteLUT[1060] = 16'hec43;
RsqrteLUT[1061] = 16'hec40;
RsqrteLUT[1062] = 16'hec3d;
RsqrteLUT[1063] = 16'hec3a;
RsqrteLUT[1064] = 16'hec38;
RsqrteLUT[1065] = 16'hec35;
RsqrteLUT[1066] = 16'hec32;
RsqrteLUT[1067] = 16'hec2f;
RsqrteLUT[1068] = 16'hec2d;
RsqrteLUT[1069] = 16'hec2a;
RsqrteLUT[1070] = 16'hec28;
RsqrteLUT[1071] = 16'hec25;
RsqrteLUT[1072] = 16'hec23;
RsqrteLUT[1073] = 16'hec20;
RsqrteLUT[1074] = 16'hec1e;
RsqrteLUT[1075] = 16'hec1c;
RsqrteLUT[1076] = 16'hec19;
RsqrteLUT[1077] = 16'hec17;
RsqrteLUT[1078] = 16'hec15;
RsqrteLUT[1079] = 16'hec13;
RsqrteLUT[1080] = 16'hec10;
RsqrteLUT[1081] = 16'hec0e;
RsqrteLUT[1082] = 16'hec0c;
RsqrteLUT[1083] = 16'hec0a;
RsqrteLUT[1084] = 16'hec08;
RsqrteLUT[1085] = 16'hec06;
RsqrteLUT[1086] = 16'hec04;
RsqrteLUT[1087] = 16'hec02;
RsqrteLUT[1088] = 16'hec00;
RsqrteLUT[1089] = 16'hebf8;
RsqrteLUT[1090] = 16'hebf0;
RsqrteLUT[1091] = 16'hebe8;
RsqrteLUT[1092] = 16'hebe1;
RsqrteLUT[1093] = 16'hebda;
RsqrteLUT[1094] = 16'hebd3;
RsqrteLUT[1095] = 16'hebcc;
RsqrteLUT[1096] = 16'hebc5;
RsqrteLUT[1097] = 16'hebbe;
RsqrteLUT[1098] = 16'hebb8;
RsqrteLUT[1099] = 16'hebb1;
RsqrteLUT[1100] = 16'hebab;
RsqrteLUT[1101] = 16'heba5;
RsqrteLUT[1102] = 16'heb9f;
RsqrteLUT[1103] = 16'heb99;
RsqrteLUT[1104] = 16'heb93;
RsqrteLUT[1105] = 16'heb8e;
RsqrteLUT[1106] = 16'heb88;
RsqrteLUT[1107] = 16'heb83;
RsqrteLUT[1108] = 16'heb7d;
RsqrteLUT[1109] = 16'heb78;
RsqrteLUT[1110] = 16'heb73;
RsqrteLUT[1111] = 16'heb6e;
RsqrteLUT[1112] = 16'heb69;
RsqrteLUT[1113] = 16'heb64;
RsqrteLUT[1114] = 16'heb5f;
RsqrteLUT[1115] = 16'heb5a;
RsqrteLUT[1116] = 16'heb56;
RsqrteLUT[1117] = 16'heb51;
RsqrteLUT[1118] = 16'heb4c;
RsqrteLUT[1119] = 16'heb48;
RsqrteLUT[1120] = 16'heb44;
RsqrteLUT[1121] = 16'heb3f;
RsqrteLUT[1122] = 16'heb3b;
RsqrteLUT[1123] = 16'heb37;
RsqrteLUT[1124] = 16'heb33;
RsqrteLUT[1125] = 16'heb2f;
RsqrteLUT[1126] = 16'heb2b;
RsqrteLUT[1127] = 16'heb27;
RsqrteLUT[1128] = 16'heb23;
RsqrteLUT[1129] = 16'heb1f;
RsqrteLUT[1130] = 16'heb1b;
RsqrteLUT[1131] = 16'heb17;
RsqrteLUT[1132] = 16'heb14;
RsqrteLUT[1133] = 16'heb10;
RsqrteLUT[1134] = 16'heb0d;
RsqrteLUT[1135] = 16'heb09;
RsqrteLUT[1136] = 16'heb06;
RsqrteLUT[1137] = 16'heb02;
RsqrteLUT[1138] = 16'heaff;
RsqrteLUT[1139] = 16'heafb;
RsqrteLUT[1140] = 16'heaf8;
RsqrteLUT[1141] = 16'heaf5;
RsqrteLUT[1142] = 16'heaf2;
RsqrteLUT[1143] = 16'heaee;
RsqrteLUT[1144] = 16'heaeb;
RsqrteLUT[1145] = 16'heae8;
RsqrteLUT[1146] = 16'heae5;
RsqrteLUT[1147] = 16'heae2;
RsqrteLUT[1148] = 16'headf;
RsqrteLUT[1149] = 16'headc;
RsqrteLUT[1150] = 16'head9;
RsqrteLUT[1151] = 16'head6;
RsqrteLUT[1152] = 16'head4;
RsqrteLUT[1153] = 16'heace;
RsqrteLUT[1154] = 16'heac9;
RsqrteLUT[1155] = 16'heac3;
RsqrteLUT[1156] = 16'heabe;
RsqrteLUT[1157] = 16'heab9;
RsqrteLUT[1158] = 16'heab4;
RsqrteLUT[1159] = 16'heaaf;
RsqrteLUT[1160] = 16'heaaa;
RsqrteLUT[1161] = 16'heaa5;
RsqrteLUT[1162] = 16'heaa1;
RsqrteLUT[1163] = 16'hea9c;
RsqrteLUT[1164] = 16'hea98;
RsqrteLUT[1165] = 16'hea94;
RsqrteLUT[1166] = 16'hea8f;
RsqrteLUT[1167] = 16'hea8b;
RsqrteLUT[1168] = 16'hea87;
RsqrteLUT[1169] = 16'hea83;
RsqrteLUT[1170] = 16'hea7f;
RsqrteLUT[1171] = 16'hea7b;
RsqrteLUT[1172] = 16'hea78;
RsqrteLUT[1173] = 16'hea74;
RsqrteLUT[1174] = 16'hea70;
RsqrteLUT[1175] = 16'hea6d;
RsqrteLUT[1176] = 16'hea69;
RsqrteLUT[1177] = 16'hea66;
RsqrteLUT[1178] = 16'hea62;
RsqrteLUT[1179] = 16'hea5f;
RsqrteLUT[1180] = 16'hea5b;
RsqrteLUT[1181] = 16'hea58;
RsqrteLUT[1182] = 16'hea55;
RsqrteLUT[1183] = 16'hea52;
RsqrteLUT[1184] = 16'hea4f;
RsqrteLUT[1185] = 16'hea4c;
RsqrteLUT[1186] = 16'hea49;
RsqrteLUT[1187] = 16'hea46;
RsqrteLUT[1188] = 16'hea43;
RsqrteLUT[1189] = 16'hea40;
RsqrteLUT[1190] = 16'hea3d;
RsqrteLUT[1191] = 16'hea3a;
RsqrteLUT[1192] = 16'hea38;
RsqrteLUT[1193] = 16'hea35;
RsqrteLUT[1194] = 16'hea32;
RsqrteLUT[1195] = 16'hea2f;
RsqrteLUT[1196] = 16'hea2d;
RsqrteLUT[1197] = 16'hea2a;
RsqrteLUT[1198] = 16'hea28;
RsqrteLUT[1199] = 16'hea25;
RsqrteLUT[1200] = 16'hea23;
RsqrteLUT[1201] = 16'hea20;
RsqrteLUT[1202] = 16'hea1e;
RsqrteLUT[1203] = 16'hea1c;
RsqrteLUT[1204] = 16'hea19;
RsqrteLUT[1205] = 16'hea17;
RsqrteLUT[1206] = 16'hea15;
RsqrteLUT[1207] = 16'hea13;
RsqrteLUT[1208] = 16'hea10;
RsqrteLUT[1209] = 16'hea0e;
RsqrteLUT[1210] = 16'hea0c;
RsqrteLUT[1211] = 16'hea0a;
RsqrteLUT[1212] = 16'hea08;
RsqrteLUT[1213] = 16'hea06;
RsqrteLUT[1214] = 16'hea04;
RsqrteLUT[1215] = 16'hea02;
RsqrteLUT[1216] = 16'hea00;
RsqrteLUT[1217] = 16'he9f8;
RsqrteLUT[1218] = 16'he9f0;
RsqrteLUT[1219] = 16'he9e8;
RsqrteLUT[1220] = 16'he9e1;
RsqrteLUT[1221] = 16'he9da;
RsqrteLUT[1222] = 16'he9d3;
RsqrteLUT[1223] = 16'he9cc;
RsqrteLUT[1224] = 16'he9c5;
RsqrteLUT[1225] = 16'he9be;
RsqrteLUT[1226] = 16'he9b8;
RsqrteLUT[1227] = 16'he9b1;
RsqrteLUT[1228] = 16'he9ab;
RsqrteLUT[1229] = 16'he9a5;
RsqrteLUT[1230] = 16'he99f;
RsqrteLUT[1231] = 16'he999;
RsqrteLUT[1232] = 16'he993;
RsqrteLUT[1233] = 16'he98e;
RsqrteLUT[1234] = 16'he988;
RsqrteLUT[1235] = 16'he983;
RsqrteLUT[1236] = 16'he97d;
RsqrteLUT[1237] = 16'he978;
RsqrteLUT[1238] = 16'he973;
RsqrteLUT[1239] = 16'he96e;
RsqrteLUT[1240] = 16'he969;
RsqrteLUT[1241] = 16'he964;
RsqrteLUT[1242] = 16'he95f;
RsqrteLUT[1243] = 16'he95a;
RsqrteLUT[1244] = 16'he956;
RsqrteLUT[1245] = 16'he951;
RsqrteLUT[1246] = 16'he94c;
RsqrteLUT[1247] = 16'he948;
RsqrteLUT[1248] = 16'he944;
RsqrteLUT[1249] = 16'he93f;
RsqrteLUT[1250] = 16'he93b;
RsqrteLUT[1251] = 16'he937;
RsqrteLUT[1252] = 16'he933;
RsqrteLUT[1253] = 16'he92f;
RsqrteLUT[1254] = 16'he92b;
RsqrteLUT[1255] = 16'he927;
RsqrteLUT[1256] = 16'he923;
RsqrteLUT[1257] = 16'he91f;
RsqrteLUT[1258] = 16'he91b;
RsqrteLUT[1259] = 16'he917;
RsqrteLUT[1260] = 16'he914;
RsqrteLUT[1261] = 16'he910;
RsqrteLUT[1262] = 16'he90d;
RsqrteLUT[1263] = 16'he909;
RsqrteLUT[1264] = 16'he906;
RsqrteLUT[1265] = 16'he902;
RsqrteLUT[1266] = 16'he8ff;
RsqrteLUT[1267] = 16'he8fb;
RsqrteLUT[1268] = 16'he8f8;
RsqrteLUT[1269] = 16'he8f5;
RsqrteLUT[1270] = 16'he8f2;
RsqrteLUT[1271] = 16'he8ee;
RsqrteLUT[1272] = 16'he8eb;
RsqrteLUT[1273] = 16'he8e8;
RsqrteLUT[1274] = 16'he8e5;
RsqrteLUT[1275] = 16'he8e2;
RsqrteLUT[1276] = 16'he8df;
RsqrteLUT[1277] = 16'he8dc;
RsqrteLUT[1278] = 16'he8d9;
RsqrteLUT[1279] = 16'he8d6;
RsqrteLUT[1280] = 16'he8d4;
RsqrteLUT[1281] = 16'he8ce;
RsqrteLUT[1282] = 16'he8c9;
RsqrteLUT[1283] = 16'he8c3;
RsqrteLUT[1284] = 16'he8be;
RsqrteLUT[1285] = 16'he8b9;
RsqrteLUT[1286] = 16'he8b4;
RsqrteLUT[1287] = 16'he8af;
RsqrteLUT[1288] = 16'he8aa;
RsqrteLUT[1289] = 16'he8a5;
RsqrteLUT[1290] = 16'he8a1;
RsqrteLUT[1291] = 16'he89c;
RsqrteLUT[1292] = 16'he898;
RsqrteLUT[1293] = 16'he894;
RsqrteLUT[1294] = 16'he88f;
RsqrteLUT[1295] = 16'he88b;
RsqrteLUT[1296] = 16'he887;
RsqrteLUT[1297] = 16'he883;
RsqrteLUT[1298] = 16'he87f;
RsqrteLUT[1299] = 16'he87b;
RsqrteLUT[1300] = 16'he878;
RsqrteLUT[1301] = 16'he874;
RsqrteLUT[1302] = 16'he870;
RsqrteLUT[1303] = 16'he86d;
RsqrteLUT[1304] = 16'he869;
RsqrteLUT[1305] = 16'he866;
RsqrteLUT[1306] = 16'he862;
RsqrteLUT[1307] = 16'he85f;
RsqrteLUT[1308] = 16'he85b;
RsqrteLUT[1309] = 16'he858;
RsqrteLUT[1310] = 16'he855;
RsqrteLUT[1311] = 16'he852;
RsqrteLUT[1312] = 16'he84f;
RsqrteLUT[1313] = 16'he84c;
RsqrteLUT[1314] = 16'he849;
RsqrteLUT[1315] = 16'he846;
RsqrteLUT[1316] = 16'he843;
RsqrteLUT[1317] = 16'he840;
RsqrteLUT[1318] = 16'he83d;
RsqrteLUT[1319] = 16'he83a;
RsqrteLUT[1320] = 16'he838;
RsqrteLUT[1321] = 16'he835;
RsqrteLUT[1322] = 16'he832;
RsqrteLUT[1323] = 16'he82f;
RsqrteLUT[1324] = 16'he82d;
RsqrteLUT[1325] = 16'he82a;
RsqrteLUT[1326] = 16'he828;
RsqrteLUT[1327] = 16'he825;
RsqrteLUT[1328] = 16'he823;
RsqrteLUT[1329] = 16'he820;
RsqrteLUT[1330] = 16'he81e;
RsqrteLUT[1331] = 16'he81c;
RsqrteLUT[1332] = 16'he819;
RsqrteLUT[1333] = 16'he817;
RsqrteLUT[1334] = 16'he815;
RsqrteLUT[1335] = 16'he813;
RsqrteLUT[1336] = 16'he810;
RsqrteLUT[1337] = 16'he80e;
RsqrteLUT[1338] = 16'he80c;
RsqrteLUT[1339] = 16'he80a;
RsqrteLUT[1340] = 16'he808;
RsqrteLUT[1341] = 16'he806;
RsqrteLUT[1342] = 16'he804;
RsqrteLUT[1343] = 16'he802;
RsqrteLUT[1344] = 16'he800;
RsqrteLUT[1345] = 16'he7f8;
RsqrteLUT[1346] = 16'he7f0;
RsqrteLUT[1347] = 16'he7e8;
RsqrteLUT[1348] = 16'he7e1;
RsqrteLUT[1349] = 16'he7da;
RsqrteLUT[1350] = 16'he7d3;
RsqrteLUT[1351] = 16'he7cc;
RsqrteLUT[1352] = 16'he7c5;
RsqrteLUT[1353] = 16'he7be;
RsqrteLUT[1354] = 16'he7b8;
RsqrteLUT[1355] = 16'he7b1;
RsqrteLUT[1356] = 16'he7ab;
RsqrteLUT[1357] = 16'he7a5;
RsqrteLUT[1358] = 16'he79f;
RsqrteLUT[1359] = 16'he799;
RsqrteLUT[1360] = 16'he793;
RsqrteLUT[1361] = 16'he78e;
RsqrteLUT[1362] = 16'he788;
RsqrteLUT[1363] = 16'he783;
RsqrteLUT[1364] = 16'he77d;
RsqrteLUT[1365] = 16'he778;
RsqrteLUT[1366] = 16'he773;
RsqrteLUT[1367] = 16'he76e;
RsqrteLUT[1368] = 16'he769;
RsqrteLUT[1369] = 16'he764;
RsqrteLUT[1370] = 16'he75f;
RsqrteLUT[1371] = 16'he75a;
RsqrteLUT[1372] = 16'he756;
RsqrteLUT[1373] = 16'he751;
RsqrteLUT[1374] = 16'he74c;
RsqrteLUT[1375] = 16'he748;
RsqrteLUT[1376] = 16'he744;
RsqrteLUT[1377] = 16'he73f;
RsqrteLUT[1378] = 16'he73b;
RsqrteLUT[1379] = 16'he737;
RsqrteLUT[1380] = 16'he733;
RsqrteLUT[1381] = 16'he72f;
RsqrteLUT[1382] = 16'he72b;
RsqrteLUT[1383] = 16'he727;
RsqrteLUT[1384] = 16'he723;
RsqrteLUT[1385] = 16'he71f;
RsqrteLUT[1386] = 16'he71b;
RsqrteLUT[1387] = 16'he717;
RsqrteLUT[1388] = 16'he714;
RsqrteLUT[1389] = 16'he710;
RsqrteLUT[1390] = 16'he70d;
RsqrteLUT[1391] = 16'he709;
RsqrteLUT[1392] = 16'he706;
RsqrteLUT[1393] = 16'he702;
RsqrteLUT[1394] = 16'he6ff;
RsqrteLUT[1395] = 16'he6fb;
RsqrteLUT[1396] = 16'he6f8;
RsqrteLUT[1397] = 16'he6f5;
RsqrteLUT[1398] = 16'he6f2;
RsqrteLUT[1399] = 16'he6ee;
RsqrteLUT[1400] = 16'he6eb;
RsqrteLUT[1401] = 16'he6e8;
RsqrteLUT[1402] = 16'he6e5;
RsqrteLUT[1403] = 16'he6e2;
RsqrteLUT[1404] = 16'he6df;
RsqrteLUT[1405] = 16'he6dc;
RsqrteLUT[1406] = 16'he6d9;
RsqrteLUT[1407] = 16'he6d6;
RsqrteLUT[1408] = 16'he6d4;
RsqrteLUT[1409] = 16'he6ce;
RsqrteLUT[1410] = 16'he6c9;
RsqrteLUT[1411] = 16'he6c3;
RsqrteLUT[1412] = 16'he6be;
RsqrteLUT[1413] = 16'he6b9;
RsqrteLUT[1414] = 16'he6b4;
RsqrteLUT[1415] = 16'he6af;
RsqrteLUT[1416] = 16'he6aa;
RsqrteLUT[1417] = 16'he6a5;
RsqrteLUT[1418] = 16'he6a1;
RsqrteLUT[1419] = 16'he69c;
RsqrteLUT[1420] = 16'he698;
RsqrteLUT[1421] = 16'he694;
RsqrteLUT[1422] = 16'he68f;
RsqrteLUT[1423] = 16'he68b;
RsqrteLUT[1424] = 16'he687;
RsqrteLUT[1425] = 16'he683;
RsqrteLUT[1426] = 16'he67f;
RsqrteLUT[1427] = 16'he67b;
RsqrteLUT[1428] = 16'he678;
RsqrteLUT[1429] = 16'he674;
RsqrteLUT[1430] = 16'he670;
RsqrteLUT[1431] = 16'he66d;
RsqrteLUT[1432] = 16'he669;
RsqrteLUT[1433] = 16'he666;
RsqrteLUT[1434] = 16'he662;
RsqrteLUT[1435] = 16'he65f;
RsqrteLUT[1436] = 16'he65b;
RsqrteLUT[1437] = 16'he658;
RsqrteLUT[1438] = 16'he655;
RsqrteLUT[1439] = 16'he652;
RsqrteLUT[1440] = 16'he64f;
RsqrteLUT[1441] = 16'he64c;
RsqrteLUT[1442] = 16'he649;
RsqrteLUT[1443] = 16'he646;
RsqrteLUT[1444] = 16'he643;
RsqrteLUT[1445] = 16'he640;
RsqrteLUT[1446] = 16'he63d;
RsqrteLUT[1447] = 16'he63a;
RsqrteLUT[1448] = 16'he638;
RsqrteLUT[1449] = 16'he635;
RsqrteLUT[1450] = 16'he632;
RsqrteLUT[1451] = 16'he62f;
RsqrteLUT[1452] = 16'he62d;
RsqrteLUT[1453] = 16'he62a;
RsqrteLUT[1454] = 16'he628;
RsqrteLUT[1455] = 16'he625;
RsqrteLUT[1456] = 16'he623;
RsqrteLUT[1457] = 16'he620;
RsqrteLUT[1458] = 16'he61e;
RsqrteLUT[1459] = 16'he61c;
RsqrteLUT[1460] = 16'he619;
RsqrteLUT[1461] = 16'he617;
RsqrteLUT[1462] = 16'he615;
RsqrteLUT[1463] = 16'he613;
RsqrteLUT[1464] = 16'he610;
RsqrteLUT[1465] = 16'he60e;
RsqrteLUT[1466] = 16'he60c;
RsqrteLUT[1467] = 16'he60a;
RsqrteLUT[1468] = 16'he608;
RsqrteLUT[1469] = 16'he606;
RsqrteLUT[1470] = 16'he604;
RsqrteLUT[1471] = 16'he602;
RsqrteLUT[1472] = 16'he600;
RsqrteLUT[1473] = 16'he5f8;
RsqrteLUT[1474] = 16'he5f0;
RsqrteLUT[1475] = 16'he5e8;
RsqrteLUT[1476] = 16'he5e1;
RsqrteLUT[1477] = 16'he5da;
RsqrteLUT[1478] = 16'he5d3;
RsqrteLUT[1479] = 16'he5cc;
RsqrteLUT[1480] = 16'he5c5;
RsqrteLUT[1481] = 16'he5be;
RsqrteLUT[1482] = 16'he5b8;
RsqrteLUT[1483] = 16'he5b1;
RsqrteLUT[1484] = 16'he5ab;
RsqrteLUT[1485] = 16'he5a5;
RsqrteLUT[1486] = 16'he59f;
RsqrteLUT[1487] = 16'he599;
RsqrteLUT[1488] = 16'he593;
RsqrteLUT[1489] = 16'he58e;
RsqrteLUT[1490] = 16'he588;
RsqrteLUT[1491] = 16'he583;
RsqrteLUT[1492] = 16'he57d;
RsqrteLUT[1493] = 16'he578;
RsqrteLUT[1494] = 16'he573;
RsqrteLUT[1495] = 16'he56e;
RsqrteLUT[1496] = 16'he569;
RsqrteLUT[1497] = 16'he564;
RsqrteLUT[1498] = 16'he55f;
RsqrteLUT[1499] = 16'he55a;
RsqrteLUT[1500] = 16'he556;
RsqrteLUT[1501] = 16'he551;
RsqrteLUT[1502] = 16'he54c;
RsqrteLUT[1503] = 16'he548;
RsqrteLUT[1504] = 16'he544;
RsqrteLUT[1505] = 16'he53f;
RsqrteLUT[1506] = 16'he53b;
RsqrteLUT[1507] = 16'he537;
RsqrteLUT[1508] = 16'he533;
RsqrteLUT[1509] = 16'he52f;
RsqrteLUT[1510] = 16'he52b;
RsqrteLUT[1511] = 16'he527;
RsqrteLUT[1512] = 16'he523;
RsqrteLUT[1513] = 16'he51f;
RsqrteLUT[1514] = 16'he51b;
RsqrteLUT[1515] = 16'he517;
RsqrteLUT[1516] = 16'he514;
RsqrteLUT[1517] = 16'he510;
RsqrteLUT[1518] = 16'he50d;
RsqrteLUT[1519] = 16'he509;
RsqrteLUT[1520] = 16'he506;
RsqrteLUT[1521] = 16'he502;
RsqrteLUT[1522] = 16'he4ff;
RsqrteLUT[1523] = 16'he4fb;
RsqrteLUT[1524] = 16'he4f8;
RsqrteLUT[1525] = 16'he4f5;
RsqrteLUT[1526] = 16'he4f2;
RsqrteLUT[1527] = 16'he4ee;
RsqrteLUT[1528] = 16'he4eb;
RsqrteLUT[1529] = 16'he4e8;
RsqrteLUT[1530] = 16'he4e5;
RsqrteLUT[1531] = 16'he4e2;
RsqrteLUT[1532] = 16'he4df;
RsqrteLUT[1533] = 16'he4dc;
RsqrteLUT[1534] = 16'he4d9;
RsqrteLUT[1535] = 16'he4d6;
RsqrteLUT[1536] = 16'he4d4;
RsqrteLUT[1537] = 16'he4ce;
RsqrteLUT[1538] = 16'he4c9;
RsqrteLUT[1539] = 16'he4c3;
RsqrteLUT[1540] = 16'he4be;
RsqrteLUT[1541] = 16'he4b9;
RsqrteLUT[1542] = 16'he4b4;
RsqrteLUT[1543] = 16'he4af;
RsqrteLUT[1544] = 16'he4aa;
RsqrteLUT[1545] = 16'he4a5;
RsqrteLUT[1546] = 16'he4a1;
RsqrteLUT[1547] = 16'he49c;
RsqrteLUT[1548] = 16'he498;
RsqrteLUT[1549] = 16'he494;
RsqrteLUT[1550] = 16'he48f;
RsqrteLUT[1551] = 16'he48b;
RsqrteLUT[1552] = 16'he487;
RsqrteLUT[1553] = 16'he483;
RsqrteLUT[1554] = 16'he47f;
RsqrteLUT[1555] = 16'he47b;
RsqrteLUT[1556] = 16'he478;
RsqrteLUT[1557] = 16'he474;
RsqrteLUT[1558] = 16'he470;
RsqrteLUT[1559] = 16'he46d;
RsqrteLUT[1560] = 16'he469;
RsqrteLUT[1561] = 16'he466;
RsqrteLUT[1562] = 16'he462;
RsqrteLUT[1563] = 16'he45f;
RsqrteLUT[1564] = 16'he45b;
RsqrteLUT[1565] = 16'he458;
RsqrteLUT[1566] = 16'he455;
RsqrteLUT[1567] = 16'he452;
RsqrteLUT[1568] = 16'he44f;
RsqrteLUT[1569] = 16'he44c;
RsqrteLUT[1570] = 16'he449;
RsqrteLUT[1571] = 16'he446;
RsqrteLUT[1572] = 16'he443;
RsqrteLUT[1573] = 16'he440;
RsqrteLUT[1574] = 16'he43d;
RsqrteLUT[1575] = 16'he43a;
RsqrteLUT[1576] = 16'he438;
RsqrteLUT[1577] = 16'he435;
RsqrteLUT[1578] = 16'he432;
RsqrteLUT[1579] = 16'he42f;
RsqrteLUT[1580] = 16'he42d;
RsqrteLUT[1581] = 16'he42a;
RsqrteLUT[1582] = 16'he428;
RsqrteLUT[1583] = 16'he425;
RsqrteLUT[1584] = 16'he423;
RsqrteLUT[1585] = 16'he420;
RsqrteLUT[1586] = 16'he41e;
RsqrteLUT[1587] = 16'he41c;
RsqrteLUT[1588] = 16'he419;
RsqrteLUT[1589] = 16'he417;
RsqrteLUT[1590] = 16'he415;
RsqrteLUT[1591] = 16'he413;
RsqrteLUT[1592] = 16'he410;
RsqrteLUT[1593] = 16'he40e;
RsqrteLUT[1594] = 16'he40c;
RsqrteLUT[1595] = 16'he40a;
RsqrteLUT[1596] = 16'he408;
RsqrteLUT[1597] = 16'he406;
RsqrteLUT[1598] = 16'he404;
RsqrteLUT[1599] = 16'he402;
RsqrteLUT[1600] = 16'he400;
RsqrteLUT[1601] = 16'he3f8;
RsqrteLUT[1602] = 16'he3f0;
RsqrteLUT[1603] = 16'he3e8;
RsqrteLUT[1604] = 16'he3e1;
RsqrteLUT[1605] = 16'he3da;
RsqrteLUT[1606] = 16'he3d3;
RsqrteLUT[1607] = 16'he3cc;
RsqrteLUT[1608] = 16'he3c5;
RsqrteLUT[1609] = 16'he3be;
RsqrteLUT[1610] = 16'he3b8;
RsqrteLUT[1611] = 16'he3b1;
RsqrteLUT[1612] = 16'he3ab;
RsqrteLUT[1613] = 16'he3a5;
RsqrteLUT[1614] = 16'he39f;
RsqrteLUT[1615] = 16'he399;
RsqrteLUT[1616] = 16'he393;
RsqrteLUT[1617] = 16'he38e;
RsqrteLUT[1618] = 16'he388;
RsqrteLUT[1619] = 16'he383;
RsqrteLUT[1620] = 16'he37d;
RsqrteLUT[1621] = 16'he378;
RsqrteLUT[1622] = 16'he373;
RsqrteLUT[1623] = 16'he36e;
RsqrteLUT[1624] = 16'he369;
RsqrteLUT[1625] = 16'he364;
RsqrteLUT[1626] = 16'he35f;
RsqrteLUT[1627] = 16'he35a;
RsqrteLUT[1628] = 16'he356;
RsqrteLUT[1629] = 16'he351;
RsqrteLUT[1630] = 16'he34c;
RsqrteLUT[1631] = 16'he348;
RsqrteLUT[1632] = 16'he344;
RsqrteLUT[1633] = 16'he33f;
RsqrteLUT[1634] = 16'he33b;
RsqrteLUT[1635] = 16'he337;
RsqrteLUT[1636] = 16'he333;
RsqrteLUT[1637] = 16'he32f;
RsqrteLUT[1638] = 16'he32b;
RsqrteLUT[1639] = 16'he327;
RsqrteLUT[1640] = 16'he323;
RsqrteLUT[1641] = 16'he31f;
RsqrteLUT[1642] = 16'he31b;
RsqrteLUT[1643] = 16'he317;
RsqrteLUT[1644] = 16'he314;
RsqrteLUT[1645] = 16'he310;
RsqrteLUT[1646] = 16'he30d;
RsqrteLUT[1647] = 16'he309;
RsqrteLUT[1648] = 16'he306;
RsqrteLUT[1649] = 16'he302;
RsqrteLUT[1650] = 16'he2ff;
RsqrteLUT[1651] = 16'he2fb;
RsqrteLUT[1652] = 16'he2f8;
RsqrteLUT[1653] = 16'he2f5;
RsqrteLUT[1654] = 16'he2f2;
RsqrteLUT[1655] = 16'he2ee;
RsqrteLUT[1656] = 16'he2eb;
RsqrteLUT[1657] = 16'he2e8;
RsqrteLUT[1658] = 16'he2e5;
RsqrteLUT[1659] = 16'he2e2;
RsqrteLUT[1660] = 16'he2df;
RsqrteLUT[1661] = 16'he2dc;
RsqrteLUT[1662] = 16'he2d9;
RsqrteLUT[1663] = 16'he2d6;
RsqrteLUT[1664] = 16'he2d4;
RsqrteLUT[1665] = 16'he2ce;
RsqrteLUT[1666] = 16'he2c9;
RsqrteLUT[1667] = 16'he2c3;
RsqrteLUT[1668] = 16'he2be;
RsqrteLUT[1669] = 16'he2b9;
RsqrteLUT[1670] = 16'he2b4;
RsqrteLUT[1671] = 16'he2af;
RsqrteLUT[1672] = 16'he2aa;
RsqrteLUT[1673] = 16'he2a5;
RsqrteLUT[1674] = 16'he2a1;
RsqrteLUT[1675] = 16'he29c;
RsqrteLUT[1676] = 16'he298;
RsqrteLUT[1677] = 16'he294;
RsqrteLUT[1678] = 16'he28f;
RsqrteLUT[1679] = 16'he28b;
RsqrteLUT[1680] = 16'he287;
RsqrteLUT[1681] = 16'he283;
RsqrteLUT[1682] = 16'he27f;
RsqrteLUT[1683] = 16'he27b;
RsqrteLUT[1684] = 16'he278;
RsqrteLUT[1685] = 16'he274;
RsqrteLUT[1686] = 16'he270;
RsqrteLUT[1687] = 16'he26d;
RsqrteLUT[1688] = 16'he269;
RsqrteLUT[1689] = 16'he266;
RsqrteLUT[1690] = 16'he262;
RsqrteLUT[1691] = 16'he25f;
RsqrteLUT[1692] = 16'he25b;
RsqrteLUT[1693] = 16'he258;
RsqrteLUT[1694] = 16'he255;
RsqrteLUT[1695] = 16'he252;
RsqrteLUT[1696] = 16'he24f;
RsqrteLUT[1697] = 16'he24c;
RsqrteLUT[1698] = 16'he249;
RsqrteLUT[1699] = 16'he246;
RsqrteLUT[1700] = 16'he243;
RsqrteLUT[1701] = 16'he240;
RsqrteLUT[1702] = 16'he23d;
RsqrteLUT[1703] = 16'he23a;
RsqrteLUT[1704] = 16'he238;
RsqrteLUT[1705] = 16'he235;
RsqrteLUT[1706] = 16'he232;
RsqrteLUT[1707] = 16'he22f;
RsqrteLUT[1708] = 16'he22d;
RsqrteLUT[1709] = 16'he22a;
RsqrteLUT[1710] = 16'he228;
RsqrteLUT[1711] = 16'he225;
RsqrteLUT[1712] = 16'he223;
RsqrteLUT[1713] = 16'he220;
RsqrteLUT[1714] = 16'he21e;
RsqrteLUT[1715] = 16'he21c;
RsqrteLUT[1716] = 16'he219;
RsqrteLUT[1717] = 16'he217;
RsqrteLUT[1718] = 16'he215;
RsqrteLUT[1719] = 16'he213;
RsqrteLUT[1720] = 16'he210;
RsqrteLUT[1721] = 16'he20e;
RsqrteLUT[1722] = 16'he20c;
RsqrteLUT[1723] = 16'he20a;
RsqrteLUT[1724] = 16'he208;
RsqrteLUT[1725] = 16'he206;
RsqrteLUT[1726] = 16'he204;
RsqrteLUT[1727] = 16'he202;
RsqrteLUT[1728] = 16'he200;
RsqrteLUT[1729] = 16'he1f8;
RsqrteLUT[1730] = 16'he1f0;
RsqrteLUT[1731] = 16'he1e8;
RsqrteLUT[1732] = 16'he1e1;
RsqrteLUT[1733] = 16'he1da;
RsqrteLUT[1734] = 16'he1d3;
RsqrteLUT[1735] = 16'he1cc;
RsqrteLUT[1736] = 16'he1c5;
RsqrteLUT[1737] = 16'he1be;
RsqrteLUT[1738] = 16'he1b8;
RsqrteLUT[1739] = 16'he1b1;
RsqrteLUT[1740] = 16'he1ab;
RsqrteLUT[1741] = 16'he1a5;
RsqrteLUT[1742] = 16'he19f;
RsqrteLUT[1743] = 16'he199;
RsqrteLUT[1744] = 16'he193;
RsqrteLUT[1745] = 16'he18e;
RsqrteLUT[1746] = 16'he188;
RsqrteLUT[1747] = 16'he183;
RsqrteLUT[1748] = 16'he17d;
RsqrteLUT[1749] = 16'he178;
RsqrteLUT[1750] = 16'he173;
RsqrteLUT[1751] = 16'he16e;
RsqrteLUT[1752] = 16'he169;
RsqrteLUT[1753] = 16'he164;
RsqrteLUT[1754] = 16'he15f;
RsqrteLUT[1755] = 16'he15a;
RsqrteLUT[1756] = 16'he156;
RsqrteLUT[1757] = 16'he151;
RsqrteLUT[1758] = 16'he14c;
RsqrteLUT[1759] = 16'he148;
RsqrteLUT[1760] = 16'he144;
RsqrteLUT[1761] = 16'he13f;
RsqrteLUT[1762] = 16'he13b;
RsqrteLUT[1763] = 16'he137;
RsqrteLUT[1764] = 16'he133;
RsqrteLUT[1765] = 16'he12f;
RsqrteLUT[1766] = 16'he12b;
RsqrteLUT[1767] = 16'he127;
RsqrteLUT[1768] = 16'he123;
RsqrteLUT[1769] = 16'he11f;
RsqrteLUT[1770] = 16'he11b;
RsqrteLUT[1771] = 16'he117;
RsqrteLUT[1772] = 16'he114;
RsqrteLUT[1773] = 16'he110;
RsqrteLUT[1774] = 16'he10d;
RsqrteLUT[1775] = 16'he109;
RsqrteLUT[1776] = 16'he106;
RsqrteLUT[1777] = 16'he102;
RsqrteLUT[1778] = 16'he0ff;
RsqrteLUT[1779] = 16'he0fb;
RsqrteLUT[1780] = 16'he0f8;
RsqrteLUT[1781] = 16'he0f5;
RsqrteLUT[1782] = 16'he0f2;
RsqrteLUT[1783] = 16'he0ee;
RsqrteLUT[1784] = 16'he0eb;
RsqrteLUT[1785] = 16'he0e8;
RsqrteLUT[1786] = 16'he0e5;
RsqrteLUT[1787] = 16'he0e2;
RsqrteLUT[1788] = 16'he0df;
RsqrteLUT[1789] = 16'he0dc;
RsqrteLUT[1790] = 16'he0d9;
RsqrteLUT[1791] = 16'he0d6;
RsqrteLUT[1792] = 16'he0d4;
RsqrteLUT[1793] = 16'he0ce;
RsqrteLUT[1794] = 16'he0c9;
RsqrteLUT[1795] = 16'he0c3;
RsqrteLUT[1796] = 16'he0be;
RsqrteLUT[1797] = 16'he0b9;
RsqrteLUT[1798] = 16'he0b4;
RsqrteLUT[1799] = 16'he0af;
RsqrteLUT[1800] = 16'he0aa;
RsqrteLUT[1801] = 16'he0a5;
RsqrteLUT[1802] = 16'he0a1;
RsqrteLUT[1803] = 16'he09c;
RsqrteLUT[1804] = 16'he098;
RsqrteLUT[1805] = 16'he094;
RsqrteLUT[1806] = 16'he08f;
RsqrteLUT[1807] = 16'he08b;
RsqrteLUT[1808] = 16'he087;
RsqrteLUT[1809] = 16'he083;
RsqrteLUT[1810] = 16'he07f;
RsqrteLUT[1811] = 16'he07b;
RsqrteLUT[1812] = 16'he078;
RsqrteLUT[1813] = 16'he074;
RsqrteLUT[1814] = 16'he070;
RsqrteLUT[1815] = 16'he06d;
RsqrteLUT[1816] = 16'he069;
RsqrteLUT[1817] = 16'he066;
RsqrteLUT[1818] = 16'he062;
RsqrteLUT[1819] = 16'he05f;
RsqrteLUT[1820] = 16'he05b;
RsqrteLUT[1821] = 16'he058;
RsqrteLUT[1822] = 16'he055;
RsqrteLUT[1823] = 16'he052;
RsqrteLUT[1824] = 16'he04f;
RsqrteLUT[1825] = 16'he04c;
RsqrteLUT[1826] = 16'he049;
RsqrteLUT[1827] = 16'he046;
RsqrteLUT[1828] = 16'he043;
RsqrteLUT[1829] = 16'he040;
RsqrteLUT[1830] = 16'he03d;
RsqrteLUT[1831] = 16'he03a;
RsqrteLUT[1832] = 16'he038;
RsqrteLUT[1833] = 16'he035;
RsqrteLUT[1834] = 16'he032;
RsqrteLUT[1835] = 16'he02f;
RsqrteLUT[1836] = 16'he02d;
RsqrteLUT[1837] = 16'he02a;
RsqrteLUT[1838] = 16'he028;
RsqrteLUT[1839] = 16'he025;
RsqrteLUT[1840] = 16'he023;
RsqrteLUT[1841] = 16'he020;
RsqrteLUT[1842] = 16'he01e;
RsqrteLUT[1843] = 16'he01c;
RsqrteLUT[1844] = 16'he019;
RsqrteLUT[1845] = 16'he017;
RsqrteLUT[1846] = 16'he015;
RsqrteLUT[1847] = 16'he013;
RsqrteLUT[1848] = 16'he010;
RsqrteLUT[1849] = 16'he00e;
RsqrteLUT[1850] = 16'he00c;
RsqrteLUT[1851] = 16'he00a;
RsqrteLUT[1852] = 16'he008;
RsqrteLUT[1853] = 16'he006;
RsqrteLUT[1854] = 16'he004;
RsqrteLUT[1855] = 16'he002;
RsqrteLUT[1856] = 16'he000;
RsqrteLUT[1857] = 16'hdff8;
RsqrteLUT[1858] = 16'hdff0;
RsqrteLUT[1859] = 16'hdfe8;
RsqrteLUT[1860] = 16'hdfe1;
RsqrteLUT[1861] = 16'hdfda;
RsqrteLUT[1862] = 16'hdfd3;
RsqrteLUT[1863] = 16'hdfcc;
RsqrteLUT[1864] = 16'hdfc5;
RsqrteLUT[1865] = 16'hdfbe;
RsqrteLUT[1866] = 16'hdfb8;
RsqrteLUT[1867] = 16'hdfb1;
RsqrteLUT[1868] = 16'hdfab;
RsqrteLUT[1869] = 16'hdfa5;
RsqrteLUT[1870] = 16'hdf9f;
RsqrteLUT[1871] = 16'hdf99;
RsqrteLUT[1872] = 16'hdf93;
RsqrteLUT[1873] = 16'hdf8e;
RsqrteLUT[1874] = 16'hdf88;
RsqrteLUT[1875] = 16'hdf83;
RsqrteLUT[1876] = 16'hdf7d;
RsqrteLUT[1877] = 16'hdf78;
RsqrteLUT[1878] = 16'hdf73;
RsqrteLUT[1879] = 16'hdf6e;
RsqrteLUT[1880] = 16'hdf69;
RsqrteLUT[1881] = 16'hdf64;
RsqrteLUT[1882] = 16'hdf5f;
RsqrteLUT[1883] = 16'hdf5a;
RsqrteLUT[1884] = 16'hdf56;
RsqrteLUT[1885] = 16'hdf51;
RsqrteLUT[1886] = 16'hdf4c;
RsqrteLUT[1887] = 16'hdf48;
RsqrteLUT[1888] = 16'hdf44;
RsqrteLUT[1889] = 16'hdf3f;
RsqrteLUT[1890] = 16'hdf3b;
RsqrteLUT[1891] = 16'hdf37;
RsqrteLUT[1892] = 16'hdf33;
RsqrteLUT[1893] = 16'hdf2f;
RsqrteLUT[1894] = 16'hdf2b;
RsqrteLUT[1895] = 16'hdf27;
RsqrteLUT[1896] = 16'hdf23;
RsqrteLUT[1897] = 16'hdf1f;
RsqrteLUT[1898] = 16'hdf1b;
RsqrteLUT[1899] = 16'hdf17;
RsqrteLUT[1900] = 16'hdf14;
RsqrteLUT[1901] = 16'hdf10;
RsqrteLUT[1902] = 16'hdf0d;
RsqrteLUT[1903] = 16'hdf09;
RsqrteLUT[1904] = 16'hdf06;
RsqrteLUT[1905] = 16'hdf02;
RsqrteLUT[1906] = 16'hdeff;
RsqrteLUT[1907] = 16'hdefb;
RsqrteLUT[1908] = 16'hdef8;
RsqrteLUT[1909] = 16'hdef5;
RsqrteLUT[1910] = 16'hdef2;
RsqrteLUT[1911] = 16'hdeee;
RsqrteLUT[1912] = 16'hdeeb;
RsqrteLUT[1913] = 16'hdee8;
RsqrteLUT[1914] = 16'hdee5;
RsqrteLUT[1915] = 16'hdee2;
RsqrteLUT[1916] = 16'hdedf;
RsqrteLUT[1917] = 16'hdedc;
RsqrteLUT[1918] = 16'hded9;
RsqrteLUT[1919] = 16'hded6;
RsqrteLUT[1920] = 16'hded4;
RsqrteLUT[1921] = 16'hdece;
RsqrteLUT[1922] = 16'hdec9;
RsqrteLUT[1923] = 16'hdec3;
RsqrteLUT[1924] = 16'hdebe;
RsqrteLUT[1925] = 16'hdeb9;
RsqrteLUT[1926] = 16'hdeb4;
RsqrteLUT[1927] = 16'hdeaf;
RsqrteLUT[1928] = 16'hdeaa;
RsqrteLUT[1929] = 16'hdea5;
RsqrteLUT[1930] = 16'hdea1;
RsqrteLUT[1931] = 16'hde9c;
RsqrteLUT[1932] = 16'hde98;
RsqrteLUT[1933] = 16'hde94;
RsqrteLUT[1934] = 16'hde8f;
RsqrteLUT[1935] = 16'hde8b;
RsqrteLUT[1936] = 16'hde87;
RsqrteLUT[1937] = 16'hde83;
RsqrteLUT[1938] = 16'hde7f;
RsqrteLUT[1939] = 16'hde7b;
RsqrteLUT[1940] = 16'hde78;
RsqrteLUT[1941] = 16'hde74;
RsqrteLUT[1942] = 16'hde70;
RsqrteLUT[1943] = 16'hde6d;
RsqrteLUT[1944] = 16'hde69;
RsqrteLUT[1945] = 16'hde66;
RsqrteLUT[1946] = 16'hde62;
RsqrteLUT[1947] = 16'hde5f;
RsqrteLUT[1948] = 16'hde5b;
RsqrteLUT[1949] = 16'hde58;
RsqrteLUT[1950] = 16'hde55;
RsqrteLUT[1951] = 16'hde52;
RsqrteLUT[1952] = 16'hde4f;
RsqrteLUT[1953] = 16'hde4c;
RsqrteLUT[1954] = 16'hde49;
RsqrteLUT[1955] = 16'hde46;
RsqrteLUT[1956] = 16'hde43;
RsqrteLUT[1957] = 16'hde40;
RsqrteLUT[1958] = 16'hde3d;
RsqrteLUT[1959] = 16'hde3a;
RsqrteLUT[1960] = 16'hde38;
RsqrteLUT[1961] = 16'hde35;
RsqrteLUT[1962] = 16'hde32;
RsqrteLUT[1963] = 16'hde2f;
RsqrteLUT[1964] = 16'hde2d;
RsqrteLUT[1965] = 16'hde2a;
RsqrteLUT[1966] = 16'hde28;
RsqrteLUT[1967] = 16'hde25;
RsqrteLUT[1968] = 16'hde23;
RsqrteLUT[1969] = 16'hde20;
RsqrteLUT[1970] = 16'hde1e;
RsqrteLUT[1971] = 16'hde1c;
RsqrteLUT[1972] = 16'hde19;
RsqrteLUT[1973] = 16'hde17;
RsqrteLUT[1974] = 16'hde15;
RsqrteLUT[1975] = 16'hde13;
RsqrteLUT[1976] = 16'hde10;
RsqrteLUT[1977] = 16'hde0e;
RsqrteLUT[1978] = 16'hde0c;
RsqrteLUT[1979] = 16'hde0a;
RsqrteLUT[1980] = 16'hde08;
RsqrteLUT[1981] = 16'hde06;
RsqrteLUT[1982] = 16'hde04;
RsqrteLUT[1983] = 16'hde02;
RsqrteLUT[1984] = 16'hde00;
RsqrteLUT[1985] = 16'hddf8;
RsqrteLUT[1986] = 16'hddf0;
RsqrteLUT[1987] = 16'hdde8;
RsqrteLUT[1988] = 16'hdde1;
RsqrteLUT[1989] = 16'hddda;
RsqrteLUT[1990] = 16'hddd3;
RsqrteLUT[1991] = 16'hddcc;
RsqrteLUT[1992] = 16'hddc5;
RsqrteLUT[1993] = 16'hddbe;
RsqrteLUT[1994] = 16'hddb8;
RsqrteLUT[1995] = 16'hddb1;
RsqrteLUT[1996] = 16'hddab;
RsqrteLUT[1997] = 16'hdda5;
RsqrteLUT[1998] = 16'hdd9f;
RsqrteLUT[1999] = 16'hdd99;
RsqrteLUT[2000] = 16'hdd93;
RsqrteLUT[2001] = 16'hdd8e;
RsqrteLUT[2002] = 16'hdd88;
RsqrteLUT[2003] = 16'hdd83;
RsqrteLUT[2004] = 16'hdd7d;
RsqrteLUT[2005] = 16'hdd78;
RsqrteLUT[2006] = 16'hdd73;
RsqrteLUT[2007] = 16'hdd6e;
RsqrteLUT[2008] = 16'hdd69;
RsqrteLUT[2009] = 16'hdd64;
RsqrteLUT[2010] = 16'hdd5f;
RsqrteLUT[2011] = 16'hdd5a;
RsqrteLUT[2012] = 16'hdd56;
RsqrteLUT[2013] = 16'hdd51;
RsqrteLUT[2014] = 16'hdd4c;
RsqrteLUT[2015] = 16'hdd48;
RsqrteLUT[2016] = 16'hdd44;
RsqrteLUT[2017] = 16'hdd3f;
RsqrteLUT[2018] = 16'hdd3b;
RsqrteLUT[2019] = 16'hdd37;
RsqrteLUT[2020] = 16'hdd33;
RsqrteLUT[2021] = 16'hdd2f;
RsqrteLUT[2022] = 16'hdd2b;
RsqrteLUT[2023] = 16'hdd27;
RsqrteLUT[2024] = 16'hdd23;
RsqrteLUT[2025] = 16'hdd1f;
RsqrteLUT[2026] = 16'hdd1b;
RsqrteLUT[2027] = 16'hdd17;
RsqrteLUT[2028] = 16'hdd14;
RsqrteLUT[2029] = 16'hdd10;
RsqrteLUT[2030] = 16'hdd0d;
RsqrteLUT[2031] = 16'hdd09;
RsqrteLUT[2032] = 16'hdd06;
RsqrteLUT[2033] = 16'hdd02;
RsqrteLUT[2034] = 16'hdcff;
RsqrteLUT[2035] = 16'hdcfb;
RsqrteLUT[2036] = 16'hdcf8;
RsqrteLUT[2037] = 16'hdcf5;
RsqrteLUT[2038] = 16'hdcf2;
RsqrteLUT[2039] = 16'hdcee;
RsqrteLUT[2040] = 16'hdceb;
RsqrteLUT[2041] = 16'hdce8;
RsqrteLUT[2042] = 16'hdce5;
RsqrteLUT[2043] = 16'hdce2;
RsqrteLUT[2044] = 16'hdcdf;
RsqrteLUT[2045] = 16'hdcdc;
RsqrteLUT[2046] = 16'hdcd9;
RsqrteLUT[2047] = 16'hdcd6;
RsqrteLUT[2048] = 16'hdcd4;
RsqrteLUT[2049] = 16'hdcce;
RsqrteLUT[2050] = 16'hdcc9;
RsqrteLUT[2051] = 16'hdcc3;
RsqrteLUT[2052] = 16'hdcbe;
RsqrteLUT[2053] = 16'hdcb9;
RsqrteLUT[2054] = 16'hdcb4;
RsqrteLUT[2055] = 16'hdcaf;
RsqrteLUT[2056] = 16'hdcaa;
RsqrteLUT[2057] = 16'hdca5;
RsqrteLUT[2058] = 16'hdca1;
RsqrteLUT[2059] = 16'hdc9c;
RsqrteLUT[2060] = 16'hdc98;
RsqrteLUT[2061] = 16'hdc94;
RsqrteLUT[2062] = 16'hdc8f;
RsqrteLUT[2063] = 16'hdc8b;
RsqrteLUT[2064] = 16'hdc87;
RsqrteLUT[2065] = 16'hdc83;
RsqrteLUT[2066] = 16'hdc7f;
RsqrteLUT[2067] = 16'hdc7b;
RsqrteLUT[2068] = 16'hdc78;
RsqrteLUT[2069] = 16'hdc74;
RsqrteLUT[2070] = 16'hdc70;
RsqrteLUT[2071] = 16'hdc6d;
RsqrteLUT[2072] = 16'hdc69;
RsqrteLUT[2073] = 16'hdc66;
RsqrteLUT[2074] = 16'hdc62;
RsqrteLUT[2075] = 16'hdc5f;
RsqrteLUT[2076] = 16'hdc5b;
RsqrteLUT[2077] = 16'hdc58;
RsqrteLUT[2078] = 16'hdc55;
RsqrteLUT[2079] = 16'hdc52;
RsqrteLUT[2080] = 16'hdc4f;
RsqrteLUT[2081] = 16'hdc4c;
RsqrteLUT[2082] = 16'hdc49;
RsqrteLUT[2083] = 16'hdc46;
RsqrteLUT[2084] = 16'hdc43;
RsqrteLUT[2085] = 16'hdc40;
RsqrteLUT[2086] = 16'hdc3d;
RsqrteLUT[2087] = 16'hdc3a;
RsqrteLUT[2088] = 16'hdc38;
RsqrteLUT[2089] = 16'hdc35;
RsqrteLUT[2090] = 16'hdc32;
RsqrteLUT[2091] = 16'hdc2f;
RsqrteLUT[2092] = 16'hdc2d;
RsqrteLUT[2093] = 16'hdc2a;
RsqrteLUT[2094] = 16'hdc28;
RsqrteLUT[2095] = 16'hdc25;
RsqrteLUT[2096] = 16'hdc23;
RsqrteLUT[2097] = 16'hdc20;
RsqrteLUT[2098] = 16'hdc1e;
RsqrteLUT[2099] = 16'hdc1c;
RsqrteLUT[2100] = 16'hdc19;
RsqrteLUT[2101] = 16'hdc17;
RsqrteLUT[2102] = 16'hdc15;
RsqrteLUT[2103] = 16'hdc13;
RsqrteLUT[2104] = 16'hdc10;
RsqrteLUT[2105] = 16'hdc0e;
RsqrteLUT[2106] = 16'hdc0c;
RsqrteLUT[2107] = 16'hdc0a;
RsqrteLUT[2108] = 16'hdc08;
RsqrteLUT[2109] = 16'hdc06;
RsqrteLUT[2110] = 16'hdc04;
RsqrteLUT[2111] = 16'hdc02;
RsqrteLUT[2112] = 16'hdc00;
RsqrteLUT[2113] = 16'hdbf8;
RsqrteLUT[2114] = 16'hdbf0;
RsqrteLUT[2115] = 16'hdbe8;
RsqrteLUT[2116] = 16'hdbe1;
RsqrteLUT[2117] = 16'hdbda;
RsqrteLUT[2118] = 16'hdbd3;
RsqrteLUT[2119] = 16'hdbcc;
RsqrteLUT[2120] = 16'hdbc5;
RsqrteLUT[2121] = 16'hdbbe;
RsqrteLUT[2122] = 16'hdbb8;
RsqrteLUT[2123] = 16'hdbb1;
RsqrteLUT[2124] = 16'hdbab;
RsqrteLUT[2125] = 16'hdba5;
RsqrteLUT[2126] = 16'hdb9f;
RsqrteLUT[2127] = 16'hdb99;
RsqrteLUT[2128] = 16'hdb93;
RsqrteLUT[2129] = 16'hdb8e;
RsqrteLUT[2130] = 16'hdb88;
RsqrteLUT[2131] = 16'hdb83;
RsqrteLUT[2132] = 16'hdb7d;
RsqrteLUT[2133] = 16'hdb78;
RsqrteLUT[2134] = 16'hdb73;
RsqrteLUT[2135] = 16'hdb6e;
RsqrteLUT[2136] = 16'hdb69;
RsqrteLUT[2137] = 16'hdb64;
RsqrteLUT[2138] = 16'hdb5f;
RsqrteLUT[2139] = 16'hdb5a;
RsqrteLUT[2140] = 16'hdb56;
RsqrteLUT[2141] = 16'hdb51;
RsqrteLUT[2142] = 16'hdb4c;
RsqrteLUT[2143] = 16'hdb48;
RsqrteLUT[2144] = 16'hdb44;
RsqrteLUT[2145] = 16'hdb3f;
RsqrteLUT[2146] = 16'hdb3b;
RsqrteLUT[2147] = 16'hdb37;
RsqrteLUT[2148] = 16'hdb33;
RsqrteLUT[2149] = 16'hdb2f;
RsqrteLUT[2150] = 16'hdb2b;
RsqrteLUT[2151] = 16'hdb27;
RsqrteLUT[2152] = 16'hdb23;
RsqrteLUT[2153] = 16'hdb1f;
RsqrteLUT[2154] = 16'hdb1b;
RsqrteLUT[2155] = 16'hdb17;
RsqrteLUT[2156] = 16'hdb14;
RsqrteLUT[2157] = 16'hdb10;
RsqrteLUT[2158] = 16'hdb0d;
RsqrteLUT[2159] = 16'hdb09;
RsqrteLUT[2160] = 16'hdb06;
RsqrteLUT[2161] = 16'hdb02;
RsqrteLUT[2162] = 16'hdaff;
RsqrteLUT[2163] = 16'hdafb;
RsqrteLUT[2164] = 16'hdaf8;
RsqrteLUT[2165] = 16'hdaf5;
RsqrteLUT[2166] = 16'hdaf2;
RsqrteLUT[2167] = 16'hdaee;
RsqrteLUT[2168] = 16'hdaeb;
RsqrteLUT[2169] = 16'hdae8;
RsqrteLUT[2170] = 16'hdae5;
RsqrteLUT[2171] = 16'hdae2;
RsqrteLUT[2172] = 16'hdadf;
RsqrteLUT[2173] = 16'hdadc;
RsqrteLUT[2174] = 16'hdad9;
RsqrteLUT[2175] = 16'hdad6;
RsqrteLUT[2176] = 16'hdad4;
RsqrteLUT[2177] = 16'hdace;
RsqrteLUT[2178] = 16'hdac9;
RsqrteLUT[2179] = 16'hdac3;
RsqrteLUT[2180] = 16'hdabe;
RsqrteLUT[2181] = 16'hdab9;
RsqrteLUT[2182] = 16'hdab4;
RsqrteLUT[2183] = 16'hdaaf;
RsqrteLUT[2184] = 16'hdaaa;
RsqrteLUT[2185] = 16'hdaa5;
RsqrteLUT[2186] = 16'hdaa1;
RsqrteLUT[2187] = 16'hda9c;
RsqrteLUT[2188] = 16'hda98;
RsqrteLUT[2189] = 16'hda94;
RsqrteLUT[2190] = 16'hda8f;
RsqrteLUT[2191] = 16'hda8b;
RsqrteLUT[2192] = 16'hda87;
RsqrteLUT[2193] = 16'hda83;
RsqrteLUT[2194] = 16'hda7f;
RsqrteLUT[2195] = 16'hda7b;
RsqrteLUT[2196] = 16'hda78;
RsqrteLUT[2197] = 16'hda74;
RsqrteLUT[2198] = 16'hda70;
RsqrteLUT[2199] = 16'hda6d;
RsqrteLUT[2200] = 16'hda69;
RsqrteLUT[2201] = 16'hda66;
RsqrteLUT[2202] = 16'hda62;
RsqrteLUT[2203] = 16'hda5f;
RsqrteLUT[2204] = 16'hda5b;
RsqrteLUT[2205] = 16'hda58;
RsqrteLUT[2206] = 16'hda55;
RsqrteLUT[2207] = 16'hda52;
RsqrteLUT[2208] = 16'hda4f;
RsqrteLUT[2209] = 16'hda4c;
RsqrteLUT[2210] = 16'hda49;
RsqrteLUT[2211] = 16'hda46;
RsqrteLUT[2212] = 16'hda43;
RsqrteLUT[2213] = 16'hda40;
RsqrteLUT[2214] = 16'hda3d;
RsqrteLUT[2215] = 16'hda3a;
RsqrteLUT[2216] = 16'hda38;
RsqrteLUT[2217] = 16'hda35;
RsqrteLUT[2218] = 16'hda32;
RsqrteLUT[2219] = 16'hda2f;
RsqrteLUT[2220] = 16'hda2d;
RsqrteLUT[2221] = 16'hda2a;
RsqrteLUT[2222] = 16'hda28;
RsqrteLUT[2223] = 16'hda25;
RsqrteLUT[2224] = 16'hda23;
RsqrteLUT[2225] = 16'hda20;
RsqrteLUT[2226] = 16'hda1e;
RsqrteLUT[2227] = 16'hda1c;
RsqrteLUT[2228] = 16'hda19;
RsqrteLUT[2229] = 16'hda17;
RsqrteLUT[2230] = 16'hda15;
RsqrteLUT[2231] = 16'hda13;
RsqrteLUT[2232] = 16'hda10;
RsqrteLUT[2233] = 16'hda0e;
RsqrteLUT[2234] = 16'hda0c;
RsqrteLUT[2235] = 16'hda0a;
RsqrteLUT[2236] = 16'hda08;
RsqrteLUT[2237] = 16'hda06;
RsqrteLUT[2238] = 16'hda04;
RsqrteLUT[2239] = 16'hda02;
RsqrteLUT[2240] = 16'hda00;
RsqrteLUT[2241] = 16'hd9f8;
RsqrteLUT[2242] = 16'hd9f0;
RsqrteLUT[2243] = 16'hd9e8;
RsqrteLUT[2244] = 16'hd9e1;
RsqrteLUT[2245] = 16'hd9da;
RsqrteLUT[2246] = 16'hd9d3;
RsqrteLUT[2247] = 16'hd9cc;
RsqrteLUT[2248] = 16'hd9c5;
RsqrteLUT[2249] = 16'hd9be;
RsqrteLUT[2250] = 16'hd9b8;
RsqrteLUT[2251] = 16'hd9b1;
RsqrteLUT[2252] = 16'hd9ab;
RsqrteLUT[2253] = 16'hd9a5;
RsqrteLUT[2254] = 16'hd99f;
RsqrteLUT[2255] = 16'hd999;
RsqrteLUT[2256] = 16'hd993;
RsqrteLUT[2257] = 16'hd98e;
RsqrteLUT[2258] = 16'hd988;
RsqrteLUT[2259] = 16'hd983;
RsqrteLUT[2260] = 16'hd97d;
RsqrteLUT[2261] = 16'hd978;
RsqrteLUT[2262] = 16'hd973;
RsqrteLUT[2263] = 16'hd96e;
RsqrteLUT[2264] = 16'hd969;
RsqrteLUT[2265] = 16'hd964;
RsqrteLUT[2266] = 16'hd95f;
RsqrteLUT[2267] = 16'hd95a;
RsqrteLUT[2268] = 16'hd956;
RsqrteLUT[2269] = 16'hd951;
RsqrteLUT[2270] = 16'hd94c;
RsqrteLUT[2271] = 16'hd948;
RsqrteLUT[2272] = 16'hd944;
RsqrteLUT[2273] = 16'hd93f;
RsqrteLUT[2274] = 16'hd93b;
RsqrteLUT[2275] = 16'hd937;
RsqrteLUT[2276] = 16'hd933;
RsqrteLUT[2277] = 16'hd92f;
RsqrteLUT[2278] = 16'hd92b;
RsqrteLUT[2279] = 16'hd927;
RsqrteLUT[2280] = 16'hd923;
RsqrteLUT[2281] = 16'hd91f;
RsqrteLUT[2282] = 16'hd91b;
RsqrteLUT[2283] = 16'hd917;
RsqrteLUT[2284] = 16'hd914;
RsqrteLUT[2285] = 16'hd910;
RsqrteLUT[2286] = 16'hd90d;
RsqrteLUT[2287] = 16'hd909;
RsqrteLUT[2288] = 16'hd906;
RsqrteLUT[2289] = 16'hd902;
RsqrteLUT[2290] = 16'hd8ff;
RsqrteLUT[2291] = 16'hd8fb;
RsqrteLUT[2292] = 16'hd8f8;
RsqrteLUT[2293] = 16'hd8f5;
RsqrteLUT[2294] = 16'hd8f2;
RsqrteLUT[2295] = 16'hd8ee;
RsqrteLUT[2296] = 16'hd8eb;
RsqrteLUT[2297] = 16'hd8e8;
RsqrteLUT[2298] = 16'hd8e5;
RsqrteLUT[2299] = 16'hd8e2;
RsqrteLUT[2300] = 16'hd8df;
RsqrteLUT[2301] = 16'hd8dc;
RsqrteLUT[2302] = 16'hd8d9;
RsqrteLUT[2303] = 16'hd8d6;
RsqrteLUT[2304] = 16'hd8d4;
RsqrteLUT[2305] = 16'hd8ce;
RsqrteLUT[2306] = 16'hd8c9;
RsqrteLUT[2307] = 16'hd8c3;
RsqrteLUT[2308] = 16'hd8be;
RsqrteLUT[2309] = 16'hd8b9;
RsqrteLUT[2310] = 16'hd8b4;
RsqrteLUT[2311] = 16'hd8af;
RsqrteLUT[2312] = 16'hd8aa;
RsqrteLUT[2313] = 16'hd8a5;
RsqrteLUT[2314] = 16'hd8a1;
RsqrteLUT[2315] = 16'hd89c;
RsqrteLUT[2316] = 16'hd898;
RsqrteLUT[2317] = 16'hd894;
RsqrteLUT[2318] = 16'hd88f;
RsqrteLUT[2319] = 16'hd88b;
RsqrteLUT[2320] = 16'hd887;
RsqrteLUT[2321] = 16'hd883;
RsqrteLUT[2322] = 16'hd87f;
RsqrteLUT[2323] = 16'hd87b;
RsqrteLUT[2324] = 16'hd878;
RsqrteLUT[2325] = 16'hd874;
RsqrteLUT[2326] = 16'hd870;
RsqrteLUT[2327] = 16'hd86d;
RsqrteLUT[2328] = 16'hd869;
RsqrteLUT[2329] = 16'hd866;
RsqrteLUT[2330] = 16'hd862;
RsqrteLUT[2331] = 16'hd85f;
RsqrteLUT[2332] = 16'hd85b;
RsqrteLUT[2333] = 16'hd858;
RsqrteLUT[2334] = 16'hd855;
RsqrteLUT[2335] = 16'hd852;
RsqrteLUT[2336] = 16'hd84f;
RsqrteLUT[2337] = 16'hd84c;
RsqrteLUT[2338] = 16'hd849;
RsqrteLUT[2339] = 16'hd846;
RsqrteLUT[2340] = 16'hd843;
RsqrteLUT[2341] = 16'hd840;
RsqrteLUT[2342] = 16'hd83d;
RsqrteLUT[2343] = 16'hd83a;
RsqrteLUT[2344] = 16'hd838;
RsqrteLUT[2345] = 16'hd835;
RsqrteLUT[2346] = 16'hd832;
RsqrteLUT[2347] = 16'hd82f;
RsqrteLUT[2348] = 16'hd82d;
RsqrteLUT[2349] = 16'hd82a;
RsqrteLUT[2350] = 16'hd828;
RsqrteLUT[2351] = 16'hd825;
RsqrteLUT[2352] = 16'hd823;
RsqrteLUT[2353] = 16'hd820;
RsqrteLUT[2354] = 16'hd81e;
RsqrteLUT[2355] = 16'hd81c;
RsqrteLUT[2356] = 16'hd819;
RsqrteLUT[2357] = 16'hd817;
RsqrteLUT[2358] = 16'hd815;
RsqrteLUT[2359] = 16'hd813;
RsqrteLUT[2360] = 16'hd810;
RsqrteLUT[2361] = 16'hd80e;
RsqrteLUT[2362] = 16'hd80c;
RsqrteLUT[2363] = 16'hd80a;
RsqrteLUT[2364] = 16'hd808;
RsqrteLUT[2365] = 16'hd806;
RsqrteLUT[2366] = 16'hd804;
RsqrteLUT[2367] = 16'hd802;
RsqrteLUT[2368] = 16'hd800;
RsqrteLUT[2369] = 16'hd7f8;
RsqrteLUT[2370] = 16'hd7f0;
RsqrteLUT[2371] = 16'hd7e8;
RsqrteLUT[2372] = 16'hd7e1;
RsqrteLUT[2373] = 16'hd7da;
RsqrteLUT[2374] = 16'hd7d3;
RsqrteLUT[2375] = 16'hd7cc;
RsqrteLUT[2376] = 16'hd7c5;
RsqrteLUT[2377] = 16'hd7be;
RsqrteLUT[2378] = 16'hd7b8;
RsqrteLUT[2379] = 16'hd7b1;
RsqrteLUT[2380] = 16'hd7ab;
RsqrteLUT[2381] = 16'hd7a5;
RsqrteLUT[2382] = 16'hd79f;
RsqrteLUT[2383] = 16'hd799;
RsqrteLUT[2384] = 16'hd793;
RsqrteLUT[2385] = 16'hd78e;
RsqrteLUT[2386] = 16'hd788;
RsqrteLUT[2387] = 16'hd783;
RsqrteLUT[2388] = 16'hd77d;
RsqrteLUT[2389] = 16'hd778;
RsqrteLUT[2390] = 16'hd773;
RsqrteLUT[2391] = 16'hd76e;
RsqrteLUT[2392] = 16'hd769;
RsqrteLUT[2393] = 16'hd764;
RsqrteLUT[2394] = 16'hd75f;
RsqrteLUT[2395] = 16'hd75a;
RsqrteLUT[2396] = 16'hd756;
RsqrteLUT[2397] = 16'hd751;
RsqrteLUT[2398] = 16'hd74c;
RsqrteLUT[2399] = 16'hd748;
RsqrteLUT[2400] = 16'hd744;
RsqrteLUT[2401] = 16'hd73f;
RsqrteLUT[2402] = 16'hd73b;
RsqrteLUT[2403] = 16'hd737;
RsqrteLUT[2404] = 16'hd733;
RsqrteLUT[2405] = 16'hd72f;
RsqrteLUT[2406] = 16'hd72b;
RsqrteLUT[2407] = 16'hd727;
RsqrteLUT[2408] = 16'hd723;
RsqrteLUT[2409] = 16'hd71f;
RsqrteLUT[2410] = 16'hd71b;
RsqrteLUT[2411] = 16'hd717;
RsqrteLUT[2412] = 16'hd714;
RsqrteLUT[2413] = 16'hd710;
RsqrteLUT[2414] = 16'hd70d;
RsqrteLUT[2415] = 16'hd709;
RsqrteLUT[2416] = 16'hd706;
RsqrteLUT[2417] = 16'hd702;
RsqrteLUT[2418] = 16'hd6ff;
RsqrteLUT[2419] = 16'hd6fb;
RsqrteLUT[2420] = 16'hd6f8;
RsqrteLUT[2421] = 16'hd6f5;
RsqrteLUT[2422] = 16'hd6f2;
RsqrteLUT[2423] = 16'hd6ee;
RsqrteLUT[2424] = 16'hd6eb;
RsqrteLUT[2425] = 16'hd6e8;
RsqrteLUT[2426] = 16'hd6e5;
RsqrteLUT[2427] = 16'hd6e2;
RsqrteLUT[2428] = 16'hd6df;
RsqrteLUT[2429] = 16'hd6dc;
RsqrteLUT[2430] = 16'hd6d9;
RsqrteLUT[2431] = 16'hd6d6;
RsqrteLUT[2432] = 16'hd6d4;
RsqrteLUT[2433] = 16'hd6ce;
RsqrteLUT[2434] = 16'hd6c9;
RsqrteLUT[2435] = 16'hd6c3;
RsqrteLUT[2436] = 16'hd6be;
RsqrteLUT[2437] = 16'hd6b9;
RsqrteLUT[2438] = 16'hd6b4;
RsqrteLUT[2439] = 16'hd6af;
RsqrteLUT[2440] = 16'hd6aa;
RsqrteLUT[2441] = 16'hd6a5;
RsqrteLUT[2442] = 16'hd6a1;
RsqrteLUT[2443] = 16'hd69c;
RsqrteLUT[2444] = 16'hd698;
RsqrteLUT[2445] = 16'hd694;
RsqrteLUT[2446] = 16'hd68f;
RsqrteLUT[2447] = 16'hd68b;
RsqrteLUT[2448] = 16'hd687;
RsqrteLUT[2449] = 16'hd683;
RsqrteLUT[2450] = 16'hd67f;
RsqrteLUT[2451] = 16'hd67b;
RsqrteLUT[2452] = 16'hd678;
RsqrteLUT[2453] = 16'hd674;
RsqrteLUT[2454] = 16'hd670;
RsqrteLUT[2455] = 16'hd66d;
RsqrteLUT[2456] = 16'hd669;
RsqrteLUT[2457] = 16'hd666;
RsqrteLUT[2458] = 16'hd662;
RsqrteLUT[2459] = 16'hd65f;
RsqrteLUT[2460] = 16'hd65b;
RsqrteLUT[2461] = 16'hd658;
RsqrteLUT[2462] = 16'hd655;
RsqrteLUT[2463] = 16'hd652;
RsqrteLUT[2464] = 16'hd64f;
RsqrteLUT[2465] = 16'hd64c;
RsqrteLUT[2466] = 16'hd649;
RsqrteLUT[2467] = 16'hd646;
RsqrteLUT[2468] = 16'hd643;
RsqrteLUT[2469] = 16'hd640;
RsqrteLUT[2470] = 16'hd63d;
RsqrteLUT[2471] = 16'hd63a;
RsqrteLUT[2472] = 16'hd638;
RsqrteLUT[2473] = 16'hd635;
RsqrteLUT[2474] = 16'hd632;
RsqrteLUT[2475] = 16'hd62f;
RsqrteLUT[2476] = 16'hd62d;
RsqrteLUT[2477] = 16'hd62a;
RsqrteLUT[2478] = 16'hd628;
RsqrteLUT[2479] = 16'hd625;
RsqrteLUT[2480] = 16'hd623;
RsqrteLUT[2481] = 16'hd620;
RsqrteLUT[2482] = 16'hd61e;
RsqrteLUT[2483] = 16'hd61c;
RsqrteLUT[2484] = 16'hd619;
RsqrteLUT[2485] = 16'hd617;
RsqrteLUT[2486] = 16'hd615;
RsqrteLUT[2487] = 16'hd613;
RsqrteLUT[2488] = 16'hd610;
RsqrteLUT[2489] = 16'hd60e;
RsqrteLUT[2490] = 16'hd60c;
RsqrteLUT[2491] = 16'hd60a;
RsqrteLUT[2492] = 16'hd608;
RsqrteLUT[2493] = 16'hd606;
RsqrteLUT[2494] = 16'hd604;
RsqrteLUT[2495] = 16'hd602;
RsqrteLUT[2496] = 16'hd600;
RsqrteLUT[2497] = 16'hd5f8;
RsqrteLUT[2498] = 16'hd5f0;
RsqrteLUT[2499] = 16'hd5e8;
RsqrteLUT[2500] = 16'hd5e1;
RsqrteLUT[2501] = 16'hd5da;
RsqrteLUT[2502] = 16'hd5d3;
RsqrteLUT[2503] = 16'hd5cc;
RsqrteLUT[2504] = 16'hd5c5;
RsqrteLUT[2505] = 16'hd5be;
RsqrteLUT[2506] = 16'hd5b8;
RsqrteLUT[2507] = 16'hd5b1;
RsqrteLUT[2508] = 16'hd5ab;
RsqrteLUT[2509] = 16'hd5a5;
RsqrteLUT[2510] = 16'hd59f;
RsqrteLUT[2511] = 16'hd599;
RsqrteLUT[2512] = 16'hd593;
RsqrteLUT[2513] = 16'hd58e;
RsqrteLUT[2514] = 16'hd588;
RsqrteLUT[2515] = 16'hd583;
RsqrteLUT[2516] = 16'hd57d;
RsqrteLUT[2517] = 16'hd578;
RsqrteLUT[2518] = 16'hd573;
RsqrteLUT[2519] = 16'hd56e;
RsqrteLUT[2520] = 16'hd569;
RsqrteLUT[2521] = 16'hd564;
RsqrteLUT[2522] = 16'hd55f;
RsqrteLUT[2523] = 16'hd55a;
RsqrteLUT[2524] = 16'hd556;
RsqrteLUT[2525] = 16'hd551;
RsqrteLUT[2526] = 16'hd54c;
RsqrteLUT[2527] = 16'hd548;
RsqrteLUT[2528] = 16'hd544;
RsqrteLUT[2529] = 16'hd53f;
RsqrteLUT[2530] = 16'hd53b;
RsqrteLUT[2531] = 16'hd537;
RsqrteLUT[2532] = 16'hd533;
RsqrteLUT[2533] = 16'hd52f;
RsqrteLUT[2534] = 16'hd52b;
RsqrteLUT[2535] = 16'hd527;
RsqrteLUT[2536] = 16'hd523;
RsqrteLUT[2537] = 16'hd51f;
RsqrteLUT[2538] = 16'hd51b;
RsqrteLUT[2539] = 16'hd517;
RsqrteLUT[2540] = 16'hd514;
RsqrteLUT[2541] = 16'hd510;
RsqrteLUT[2542] = 16'hd50d;
RsqrteLUT[2543] = 16'hd509;
RsqrteLUT[2544] = 16'hd506;
RsqrteLUT[2545] = 16'hd502;
RsqrteLUT[2546] = 16'hd4ff;
RsqrteLUT[2547] = 16'hd4fb;
RsqrteLUT[2548] = 16'hd4f8;
RsqrteLUT[2549] = 16'hd4f5;
RsqrteLUT[2550] = 16'hd4f2;
RsqrteLUT[2551] = 16'hd4ee;
RsqrteLUT[2552] = 16'hd4eb;
RsqrteLUT[2553] = 16'hd4e8;
RsqrteLUT[2554] = 16'hd4e5;
RsqrteLUT[2555] = 16'hd4e2;
RsqrteLUT[2556] = 16'hd4df;
RsqrteLUT[2557] = 16'hd4dc;
RsqrteLUT[2558] = 16'hd4d9;
RsqrteLUT[2559] = 16'hd4d6;
RsqrteLUT[2560] = 16'hd4d4;
RsqrteLUT[2561] = 16'hd4ce;
RsqrteLUT[2562] = 16'hd4c9;
RsqrteLUT[2563] = 16'hd4c3;
RsqrteLUT[2564] = 16'hd4be;
RsqrteLUT[2565] = 16'hd4b9;
RsqrteLUT[2566] = 16'hd4b4;
RsqrteLUT[2567] = 16'hd4af;
RsqrteLUT[2568] = 16'hd4aa;
RsqrteLUT[2569] = 16'hd4a5;
RsqrteLUT[2570] = 16'hd4a1;
RsqrteLUT[2571] = 16'hd49c;
RsqrteLUT[2572] = 16'hd498;
RsqrteLUT[2573] = 16'hd494;
RsqrteLUT[2574] = 16'hd48f;
RsqrteLUT[2575] = 16'hd48b;
RsqrteLUT[2576] = 16'hd487;
RsqrteLUT[2577] = 16'hd483;
RsqrteLUT[2578] = 16'hd47f;
RsqrteLUT[2579] = 16'hd47b;
RsqrteLUT[2580] = 16'hd478;
RsqrteLUT[2581] = 16'hd474;
RsqrteLUT[2582] = 16'hd470;
RsqrteLUT[2583] = 16'hd46d;
RsqrteLUT[2584] = 16'hd469;
RsqrteLUT[2585] = 16'hd466;
RsqrteLUT[2586] = 16'hd462;
RsqrteLUT[2587] = 16'hd45f;
RsqrteLUT[2588] = 16'hd45b;
RsqrteLUT[2589] = 16'hd458;
RsqrteLUT[2590] = 16'hd455;
RsqrteLUT[2591] = 16'hd452;
RsqrteLUT[2592] = 16'hd44f;
RsqrteLUT[2593] = 16'hd44c;
RsqrteLUT[2594] = 16'hd449;
RsqrteLUT[2595] = 16'hd446;
RsqrteLUT[2596] = 16'hd443;
RsqrteLUT[2597] = 16'hd440;
RsqrteLUT[2598] = 16'hd43d;
RsqrteLUT[2599] = 16'hd43a;
RsqrteLUT[2600] = 16'hd438;
RsqrteLUT[2601] = 16'hd435;
RsqrteLUT[2602] = 16'hd432;
RsqrteLUT[2603] = 16'hd42f;
RsqrteLUT[2604] = 16'hd42d;
RsqrteLUT[2605] = 16'hd42a;
RsqrteLUT[2606] = 16'hd428;
RsqrteLUT[2607] = 16'hd425;
RsqrteLUT[2608] = 16'hd423;
RsqrteLUT[2609] = 16'hd420;
RsqrteLUT[2610] = 16'hd41e;
RsqrteLUT[2611] = 16'hd41c;
RsqrteLUT[2612] = 16'hd419;
RsqrteLUT[2613] = 16'hd417;
RsqrteLUT[2614] = 16'hd415;
RsqrteLUT[2615] = 16'hd413;
RsqrteLUT[2616] = 16'hd410;
RsqrteLUT[2617] = 16'hd40e;
RsqrteLUT[2618] = 16'hd40c;
RsqrteLUT[2619] = 16'hd40a;
RsqrteLUT[2620] = 16'hd408;
RsqrteLUT[2621] = 16'hd406;
RsqrteLUT[2622] = 16'hd404;
RsqrteLUT[2623] = 16'hd402;
RsqrteLUT[2624] = 16'hd400;
RsqrteLUT[2625] = 16'hd3f8;
RsqrteLUT[2626] = 16'hd3f0;
RsqrteLUT[2627] = 16'hd3e8;
RsqrteLUT[2628] = 16'hd3e1;
RsqrteLUT[2629] = 16'hd3da;
RsqrteLUT[2630] = 16'hd3d3;
RsqrteLUT[2631] = 16'hd3cc;
RsqrteLUT[2632] = 16'hd3c5;
RsqrteLUT[2633] = 16'hd3be;
RsqrteLUT[2634] = 16'hd3b8;
RsqrteLUT[2635] = 16'hd3b1;
RsqrteLUT[2636] = 16'hd3ab;
RsqrteLUT[2637] = 16'hd3a5;
RsqrteLUT[2638] = 16'hd39f;
RsqrteLUT[2639] = 16'hd399;
RsqrteLUT[2640] = 16'hd393;
RsqrteLUT[2641] = 16'hd38e;
RsqrteLUT[2642] = 16'hd388;
RsqrteLUT[2643] = 16'hd383;
RsqrteLUT[2644] = 16'hd37d;
RsqrteLUT[2645] = 16'hd378;
RsqrteLUT[2646] = 16'hd373;
RsqrteLUT[2647] = 16'hd36e;
RsqrteLUT[2648] = 16'hd369;
RsqrteLUT[2649] = 16'hd364;
RsqrteLUT[2650] = 16'hd35f;
RsqrteLUT[2651] = 16'hd35a;
RsqrteLUT[2652] = 16'hd356;
RsqrteLUT[2653] = 16'hd351;
RsqrteLUT[2654] = 16'hd34c;
RsqrteLUT[2655] = 16'hd348;
RsqrteLUT[2656] = 16'hd344;
RsqrteLUT[2657] = 16'hd33f;
RsqrteLUT[2658] = 16'hd33b;
RsqrteLUT[2659] = 16'hd337;
RsqrteLUT[2660] = 16'hd333;
RsqrteLUT[2661] = 16'hd32f;
RsqrteLUT[2662] = 16'hd32b;
RsqrteLUT[2663] = 16'hd327;
RsqrteLUT[2664] = 16'hd323;
RsqrteLUT[2665] = 16'hd31f;
RsqrteLUT[2666] = 16'hd31b;
RsqrteLUT[2667] = 16'hd317;
RsqrteLUT[2668] = 16'hd314;
RsqrteLUT[2669] = 16'hd310;
RsqrteLUT[2670] = 16'hd30d;
RsqrteLUT[2671] = 16'hd309;
RsqrteLUT[2672] = 16'hd306;
RsqrteLUT[2673] = 16'hd302;
RsqrteLUT[2674] = 16'hd2ff;
RsqrteLUT[2675] = 16'hd2fb;
RsqrteLUT[2676] = 16'hd2f8;
RsqrteLUT[2677] = 16'hd2f5;
RsqrteLUT[2678] = 16'hd2f2;
RsqrteLUT[2679] = 16'hd2ee;
RsqrteLUT[2680] = 16'hd2eb;
RsqrteLUT[2681] = 16'hd2e8;
RsqrteLUT[2682] = 16'hd2e5;
RsqrteLUT[2683] = 16'hd2e2;
RsqrteLUT[2684] = 16'hd2df;
RsqrteLUT[2685] = 16'hd2dc;
RsqrteLUT[2686] = 16'hd2d9;
RsqrteLUT[2687] = 16'hd2d6;
RsqrteLUT[2688] = 16'hd2d4;
RsqrteLUT[2689] = 16'hd2ce;
RsqrteLUT[2690] = 16'hd2c9;
RsqrteLUT[2691] = 16'hd2c3;
RsqrteLUT[2692] = 16'hd2be;
RsqrteLUT[2693] = 16'hd2b9;
RsqrteLUT[2694] = 16'hd2b4;
RsqrteLUT[2695] = 16'hd2af;
RsqrteLUT[2696] = 16'hd2aa;
RsqrteLUT[2697] = 16'hd2a5;
RsqrteLUT[2698] = 16'hd2a1;
RsqrteLUT[2699] = 16'hd29c;
RsqrteLUT[2700] = 16'hd298;
RsqrteLUT[2701] = 16'hd294;
RsqrteLUT[2702] = 16'hd28f;
RsqrteLUT[2703] = 16'hd28b;
RsqrteLUT[2704] = 16'hd287;
RsqrteLUT[2705] = 16'hd283;
RsqrteLUT[2706] = 16'hd27f;
RsqrteLUT[2707] = 16'hd27b;
RsqrteLUT[2708] = 16'hd278;
RsqrteLUT[2709] = 16'hd274;
RsqrteLUT[2710] = 16'hd270;
RsqrteLUT[2711] = 16'hd26d;
RsqrteLUT[2712] = 16'hd269;
RsqrteLUT[2713] = 16'hd266;
RsqrteLUT[2714] = 16'hd262;
RsqrteLUT[2715] = 16'hd25f;
RsqrteLUT[2716] = 16'hd25b;
RsqrteLUT[2717] = 16'hd258;
RsqrteLUT[2718] = 16'hd255;
RsqrteLUT[2719] = 16'hd252;
RsqrteLUT[2720] = 16'hd24f;
RsqrteLUT[2721] = 16'hd24c;
RsqrteLUT[2722] = 16'hd249;
RsqrteLUT[2723] = 16'hd246;
RsqrteLUT[2724] = 16'hd243;
RsqrteLUT[2725] = 16'hd240;
RsqrteLUT[2726] = 16'hd23d;
RsqrteLUT[2727] = 16'hd23a;
RsqrteLUT[2728] = 16'hd238;
RsqrteLUT[2729] = 16'hd235;
RsqrteLUT[2730] = 16'hd232;
RsqrteLUT[2731] = 16'hd22f;
RsqrteLUT[2732] = 16'hd22d;
RsqrteLUT[2733] = 16'hd22a;
RsqrteLUT[2734] = 16'hd228;
RsqrteLUT[2735] = 16'hd225;
RsqrteLUT[2736] = 16'hd223;
RsqrteLUT[2737] = 16'hd220;
RsqrteLUT[2738] = 16'hd21e;
RsqrteLUT[2739] = 16'hd21c;
RsqrteLUT[2740] = 16'hd219;
RsqrteLUT[2741] = 16'hd217;
RsqrteLUT[2742] = 16'hd215;
RsqrteLUT[2743] = 16'hd213;
RsqrteLUT[2744] = 16'hd210;
RsqrteLUT[2745] = 16'hd20e;
RsqrteLUT[2746] = 16'hd20c;
RsqrteLUT[2747] = 16'hd20a;
RsqrteLUT[2748] = 16'hd208;
RsqrteLUT[2749] = 16'hd206;
RsqrteLUT[2750] = 16'hd204;
RsqrteLUT[2751] = 16'hd202;
RsqrteLUT[2752] = 16'hd200;
RsqrteLUT[2753] = 16'hd1f8;
RsqrteLUT[2754] = 16'hd1f0;
RsqrteLUT[2755] = 16'hd1e8;
RsqrteLUT[2756] = 16'hd1e1;
RsqrteLUT[2757] = 16'hd1da;
RsqrteLUT[2758] = 16'hd1d3;
RsqrteLUT[2759] = 16'hd1cc;
RsqrteLUT[2760] = 16'hd1c5;
RsqrteLUT[2761] = 16'hd1be;
RsqrteLUT[2762] = 16'hd1b8;
RsqrteLUT[2763] = 16'hd1b1;
RsqrteLUT[2764] = 16'hd1ab;
RsqrteLUT[2765] = 16'hd1a5;
RsqrteLUT[2766] = 16'hd19f;
RsqrteLUT[2767] = 16'hd199;
RsqrteLUT[2768] = 16'hd193;
RsqrteLUT[2769] = 16'hd18e;
RsqrteLUT[2770] = 16'hd188;
RsqrteLUT[2771] = 16'hd183;
RsqrteLUT[2772] = 16'hd17d;
RsqrteLUT[2773] = 16'hd178;
RsqrteLUT[2774] = 16'hd173;
RsqrteLUT[2775] = 16'hd16e;
RsqrteLUT[2776] = 16'hd169;
RsqrteLUT[2777] = 16'hd164;
RsqrteLUT[2778] = 16'hd15f;
RsqrteLUT[2779] = 16'hd15a;
RsqrteLUT[2780] = 16'hd156;
RsqrteLUT[2781] = 16'hd151;
RsqrteLUT[2782] = 16'hd14c;
RsqrteLUT[2783] = 16'hd148;
RsqrteLUT[2784] = 16'hd144;
RsqrteLUT[2785] = 16'hd13f;
RsqrteLUT[2786] = 16'hd13b;
RsqrteLUT[2787] = 16'hd137;
RsqrteLUT[2788] = 16'hd133;
RsqrteLUT[2789] = 16'hd12f;
RsqrteLUT[2790] = 16'hd12b;
RsqrteLUT[2791] = 16'hd127;
RsqrteLUT[2792] = 16'hd123;
RsqrteLUT[2793] = 16'hd11f;
RsqrteLUT[2794] = 16'hd11b;
RsqrteLUT[2795] = 16'hd117;
RsqrteLUT[2796] = 16'hd114;
RsqrteLUT[2797] = 16'hd110;
RsqrteLUT[2798] = 16'hd10d;
RsqrteLUT[2799] = 16'hd109;
RsqrteLUT[2800] = 16'hd106;
RsqrteLUT[2801] = 16'hd102;
RsqrteLUT[2802] = 16'hd0ff;
RsqrteLUT[2803] = 16'hd0fb;
RsqrteLUT[2804] = 16'hd0f8;
RsqrteLUT[2805] = 16'hd0f5;
RsqrteLUT[2806] = 16'hd0f2;
RsqrteLUT[2807] = 16'hd0ee;
RsqrteLUT[2808] = 16'hd0eb;
RsqrteLUT[2809] = 16'hd0e8;
RsqrteLUT[2810] = 16'hd0e5;
RsqrteLUT[2811] = 16'hd0e2;
RsqrteLUT[2812] = 16'hd0df;
RsqrteLUT[2813] = 16'hd0dc;
RsqrteLUT[2814] = 16'hd0d9;
RsqrteLUT[2815] = 16'hd0d6;
RsqrteLUT[2816] = 16'hd0d4;
RsqrteLUT[2817] = 16'hd0ce;
RsqrteLUT[2818] = 16'hd0c9;
RsqrteLUT[2819] = 16'hd0c3;
RsqrteLUT[2820] = 16'hd0be;
RsqrteLUT[2821] = 16'hd0b9;
RsqrteLUT[2822] = 16'hd0b4;
RsqrteLUT[2823] = 16'hd0af;
RsqrteLUT[2824] = 16'hd0aa;
RsqrteLUT[2825] = 16'hd0a5;
RsqrteLUT[2826] = 16'hd0a1;
RsqrteLUT[2827] = 16'hd09c;
RsqrteLUT[2828] = 16'hd098;
RsqrteLUT[2829] = 16'hd094;
RsqrteLUT[2830] = 16'hd08f;
RsqrteLUT[2831] = 16'hd08b;
RsqrteLUT[2832] = 16'hd087;
RsqrteLUT[2833] = 16'hd083;
RsqrteLUT[2834] = 16'hd07f;
RsqrteLUT[2835] = 16'hd07b;
RsqrteLUT[2836] = 16'hd078;
RsqrteLUT[2837] = 16'hd074;
RsqrteLUT[2838] = 16'hd070;
RsqrteLUT[2839] = 16'hd06d;
RsqrteLUT[2840] = 16'hd069;
RsqrteLUT[2841] = 16'hd066;
RsqrteLUT[2842] = 16'hd062;
RsqrteLUT[2843] = 16'hd05f;
RsqrteLUT[2844] = 16'hd05b;
RsqrteLUT[2845] = 16'hd058;
RsqrteLUT[2846] = 16'hd055;
RsqrteLUT[2847] = 16'hd052;
RsqrteLUT[2848] = 16'hd04f;
RsqrteLUT[2849] = 16'hd04c;
RsqrteLUT[2850] = 16'hd049;
RsqrteLUT[2851] = 16'hd046;
RsqrteLUT[2852] = 16'hd043;
RsqrteLUT[2853] = 16'hd040;
RsqrteLUT[2854] = 16'hd03d;
RsqrteLUT[2855] = 16'hd03a;
RsqrteLUT[2856] = 16'hd038;
RsqrteLUT[2857] = 16'hd035;
RsqrteLUT[2858] = 16'hd032;
RsqrteLUT[2859] = 16'hd02f;
RsqrteLUT[2860] = 16'hd02d;
RsqrteLUT[2861] = 16'hd02a;
RsqrteLUT[2862] = 16'hd028;
RsqrteLUT[2863] = 16'hd025;
RsqrteLUT[2864] = 16'hd023;
RsqrteLUT[2865] = 16'hd020;
RsqrteLUT[2866] = 16'hd01e;
RsqrteLUT[2867] = 16'hd01c;
RsqrteLUT[2868] = 16'hd019;
RsqrteLUT[2869] = 16'hd017;
RsqrteLUT[2870] = 16'hd015;
RsqrteLUT[2871] = 16'hd013;
RsqrteLUT[2872] = 16'hd010;
RsqrteLUT[2873] = 16'hd00e;
RsqrteLUT[2874] = 16'hd00c;
RsqrteLUT[2875] = 16'hd00a;
RsqrteLUT[2876] = 16'hd008;
RsqrteLUT[2877] = 16'hd006;
RsqrteLUT[2878] = 16'hd004;
RsqrteLUT[2879] = 16'hd002;
RsqrteLUT[2880] = 16'hd000;
RsqrteLUT[2881] = 16'hcff8;
RsqrteLUT[2882] = 16'hcff0;
RsqrteLUT[2883] = 16'hcfe8;
RsqrteLUT[2884] = 16'hcfe1;
RsqrteLUT[2885] = 16'hcfda;
RsqrteLUT[2886] = 16'hcfd3;
RsqrteLUT[2887] = 16'hcfcc;
RsqrteLUT[2888] = 16'hcfc5;
RsqrteLUT[2889] = 16'hcfbe;
RsqrteLUT[2890] = 16'hcfb8;
RsqrteLUT[2891] = 16'hcfb1;
RsqrteLUT[2892] = 16'hcfab;
RsqrteLUT[2893] = 16'hcfa5;
RsqrteLUT[2894] = 16'hcf9f;
RsqrteLUT[2895] = 16'hcf99;
RsqrteLUT[2896] = 16'hcf93;
RsqrteLUT[2897] = 16'hcf8e;
RsqrteLUT[2898] = 16'hcf88;
RsqrteLUT[2899] = 16'hcf83;
RsqrteLUT[2900] = 16'hcf7d;
RsqrteLUT[2901] = 16'hcf78;
RsqrteLUT[2902] = 16'hcf73;
RsqrteLUT[2903] = 16'hcf6e;
RsqrteLUT[2904] = 16'hcf69;
RsqrteLUT[2905] = 16'hcf64;
RsqrteLUT[2906] = 16'hcf5f;
RsqrteLUT[2907] = 16'hcf5a;
RsqrteLUT[2908] = 16'hcf56;
RsqrteLUT[2909] = 16'hcf51;
RsqrteLUT[2910] = 16'hcf4c;
RsqrteLUT[2911] = 16'hcf48;
RsqrteLUT[2912] = 16'hcf44;
RsqrteLUT[2913] = 16'hcf3f;
RsqrteLUT[2914] = 16'hcf3b;
RsqrteLUT[2915] = 16'hcf37;
RsqrteLUT[2916] = 16'hcf33;
RsqrteLUT[2917] = 16'hcf2f;
RsqrteLUT[2918] = 16'hcf2b;
RsqrteLUT[2919] = 16'hcf27;
RsqrteLUT[2920] = 16'hcf23;
RsqrteLUT[2921] = 16'hcf1f;
RsqrteLUT[2922] = 16'hcf1b;
RsqrteLUT[2923] = 16'hcf17;
RsqrteLUT[2924] = 16'hcf14;
RsqrteLUT[2925] = 16'hcf10;
RsqrteLUT[2926] = 16'hcf0d;
RsqrteLUT[2927] = 16'hcf09;
RsqrteLUT[2928] = 16'hcf06;
RsqrteLUT[2929] = 16'hcf02;
RsqrteLUT[2930] = 16'hceff;
RsqrteLUT[2931] = 16'hcefb;
RsqrteLUT[2932] = 16'hcef8;
RsqrteLUT[2933] = 16'hcef5;
RsqrteLUT[2934] = 16'hcef2;
RsqrteLUT[2935] = 16'hceee;
RsqrteLUT[2936] = 16'hceeb;
RsqrteLUT[2937] = 16'hcee8;
RsqrteLUT[2938] = 16'hcee5;
RsqrteLUT[2939] = 16'hcee2;
RsqrteLUT[2940] = 16'hcedf;
RsqrteLUT[2941] = 16'hcedc;
RsqrteLUT[2942] = 16'hced9;
RsqrteLUT[2943] = 16'hced6;
RsqrteLUT[2944] = 16'hced4;
RsqrteLUT[2945] = 16'hcece;
RsqrteLUT[2946] = 16'hcec9;
RsqrteLUT[2947] = 16'hcec3;
RsqrteLUT[2948] = 16'hcebe;
RsqrteLUT[2949] = 16'hceb9;
RsqrteLUT[2950] = 16'hceb4;
RsqrteLUT[2951] = 16'hceaf;
RsqrteLUT[2952] = 16'hceaa;
RsqrteLUT[2953] = 16'hcea5;
RsqrteLUT[2954] = 16'hcea1;
RsqrteLUT[2955] = 16'hce9c;
RsqrteLUT[2956] = 16'hce98;
RsqrteLUT[2957] = 16'hce94;
RsqrteLUT[2958] = 16'hce8f;
RsqrteLUT[2959] = 16'hce8b;
RsqrteLUT[2960] = 16'hce87;
RsqrteLUT[2961] = 16'hce83;
RsqrteLUT[2962] = 16'hce7f;
RsqrteLUT[2963] = 16'hce7b;
RsqrteLUT[2964] = 16'hce78;
RsqrteLUT[2965] = 16'hce74;
RsqrteLUT[2966] = 16'hce70;
RsqrteLUT[2967] = 16'hce6d;
RsqrteLUT[2968] = 16'hce69;
RsqrteLUT[2969] = 16'hce66;
RsqrteLUT[2970] = 16'hce62;
RsqrteLUT[2971] = 16'hce5f;
RsqrteLUT[2972] = 16'hce5b;
RsqrteLUT[2973] = 16'hce58;
RsqrteLUT[2974] = 16'hce55;
RsqrteLUT[2975] = 16'hce52;
RsqrteLUT[2976] = 16'hce4f;
RsqrteLUT[2977] = 16'hce4c;
RsqrteLUT[2978] = 16'hce49;
RsqrteLUT[2979] = 16'hce46;
RsqrteLUT[2980] = 16'hce43;
RsqrteLUT[2981] = 16'hce40;
RsqrteLUT[2982] = 16'hce3d;
RsqrteLUT[2983] = 16'hce3a;
RsqrteLUT[2984] = 16'hce38;
RsqrteLUT[2985] = 16'hce35;
RsqrteLUT[2986] = 16'hce32;
RsqrteLUT[2987] = 16'hce2f;
RsqrteLUT[2988] = 16'hce2d;
RsqrteLUT[2989] = 16'hce2a;
RsqrteLUT[2990] = 16'hce28;
RsqrteLUT[2991] = 16'hce25;
RsqrteLUT[2992] = 16'hce23;
RsqrteLUT[2993] = 16'hce20;
RsqrteLUT[2994] = 16'hce1e;
RsqrteLUT[2995] = 16'hce1c;
RsqrteLUT[2996] = 16'hce19;
RsqrteLUT[2997] = 16'hce17;
RsqrteLUT[2998] = 16'hce15;
RsqrteLUT[2999] = 16'hce13;
RsqrteLUT[3000] = 16'hce10;
RsqrteLUT[3001] = 16'hce0e;
RsqrteLUT[3002] = 16'hce0c;
RsqrteLUT[3003] = 16'hce0a;
RsqrteLUT[3004] = 16'hce08;
RsqrteLUT[3005] = 16'hce06;
RsqrteLUT[3006] = 16'hce04;
RsqrteLUT[3007] = 16'hce02;
RsqrteLUT[3008] = 16'hce00;
RsqrteLUT[3009] = 16'hcdf8;
RsqrteLUT[3010] = 16'hcdf0;
RsqrteLUT[3011] = 16'hcde8;
RsqrteLUT[3012] = 16'hcde1;
RsqrteLUT[3013] = 16'hcdda;
RsqrteLUT[3014] = 16'hcdd3;
RsqrteLUT[3015] = 16'hcdcc;
RsqrteLUT[3016] = 16'hcdc5;
RsqrteLUT[3017] = 16'hcdbe;
RsqrteLUT[3018] = 16'hcdb8;
RsqrteLUT[3019] = 16'hcdb1;
RsqrteLUT[3020] = 16'hcdab;
RsqrteLUT[3021] = 16'hcda5;
RsqrteLUT[3022] = 16'hcd9f;
RsqrteLUT[3023] = 16'hcd99;
RsqrteLUT[3024] = 16'hcd93;
RsqrteLUT[3025] = 16'hcd8e;
RsqrteLUT[3026] = 16'hcd88;
RsqrteLUT[3027] = 16'hcd83;
RsqrteLUT[3028] = 16'hcd7d;
RsqrteLUT[3029] = 16'hcd78;
RsqrteLUT[3030] = 16'hcd73;
RsqrteLUT[3031] = 16'hcd6e;
RsqrteLUT[3032] = 16'hcd69;
RsqrteLUT[3033] = 16'hcd64;
RsqrteLUT[3034] = 16'hcd5f;
RsqrteLUT[3035] = 16'hcd5a;
RsqrteLUT[3036] = 16'hcd56;
RsqrteLUT[3037] = 16'hcd51;
RsqrteLUT[3038] = 16'hcd4c;
RsqrteLUT[3039] = 16'hcd48;
RsqrteLUT[3040] = 16'hcd44;
RsqrteLUT[3041] = 16'hcd3f;
RsqrteLUT[3042] = 16'hcd3b;
RsqrteLUT[3043] = 16'hcd37;
RsqrteLUT[3044] = 16'hcd33;
RsqrteLUT[3045] = 16'hcd2f;
RsqrteLUT[3046] = 16'hcd2b;
RsqrteLUT[3047] = 16'hcd27;
RsqrteLUT[3048] = 16'hcd23;
RsqrteLUT[3049] = 16'hcd1f;
RsqrteLUT[3050] = 16'hcd1b;
RsqrteLUT[3051] = 16'hcd17;
RsqrteLUT[3052] = 16'hcd14;
RsqrteLUT[3053] = 16'hcd10;
RsqrteLUT[3054] = 16'hcd0d;
RsqrteLUT[3055] = 16'hcd09;
RsqrteLUT[3056] = 16'hcd06;
RsqrteLUT[3057] = 16'hcd02;
RsqrteLUT[3058] = 16'hccff;
RsqrteLUT[3059] = 16'hccfb;
RsqrteLUT[3060] = 16'hccf8;
RsqrteLUT[3061] = 16'hccf5;
RsqrteLUT[3062] = 16'hccf2;
RsqrteLUT[3063] = 16'hccee;
RsqrteLUT[3064] = 16'hcceb;
RsqrteLUT[3065] = 16'hcce8;
RsqrteLUT[3066] = 16'hcce5;
RsqrteLUT[3067] = 16'hcce2;
RsqrteLUT[3068] = 16'hccdf;
RsqrteLUT[3069] = 16'hccdc;
RsqrteLUT[3070] = 16'hccd9;
RsqrteLUT[3071] = 16'hccd6;
RsqrteLUT[3072] = 16'hccd4;
RsqrteLUT[3073] = 16'hccce;
RsqrteLUT[3074] = 16'hccc9;
RsqrteLUT[3075] = 16'hccc3;
RsqrteLUT[3076] = 16'hccbe;
RsqrteLUT[3077] = 16'hccb9;
RsqrteLUT[3078] = 16'hccb4;
RsqrteLUT[3079] = 16'hccaf;
RsqrteLUT[3080] = 16'hccaa;
RsqrteLUT[3081] = 16'hcca5;
RsqrteLUT[3082] = 16'hcca1;
RsqrteLUT[3083] = 16'hcc9c;
RsqrteLUT[3084] = 16'hcc98;
RsqrteLUT[3085] = 16'hcc94;
RsqrteLUT[3086] = 16'hcc8f;
RsqrteLUT[3087] = 16'hcc8b;
RsqrteLUT[3088] = 16'hcc87;
RsqrteLUT[3089] = 16'hcc83;
RsqrteLUT[3090] = 16'hcc7f;
RsqrteLUT[3091] = 16'hcc7b;
RsqrteLUT[3092] = 16'hcc78;
RsqrteLUT[3093] = 16'hcc74;
RsqrteLUT[3094] = 16'hcc70;
RsqrteLUT[3095] = 16'hcc6d;
RsqrteLUT[3096] = 16'hcc69;
RsqrteLUT[3097] = 16'hcc66;
RsqrteLUT[3098] = 16'hcc62;
RsqrteLUT[3099] = 16'hcc5f;
RsqrteLUT[3100] = 16'hcc5b;
RsqrteLUT[3101] = 16'hcc58;
RsqrteLUT[3102] = 16'hcc55;
RsqrteLUT[3103] = 16'hcc52;
RsqrteLUT[3104] = 16'hcc4f;
RsqrteLUT[3105] = 16'hcc4c;
RsqrteLUT[3106] = 16'hcc49;
RsqrteLUT[3107] = 16'hcc46;
RsqrteLUT[3108] = 16'hcc43;
RsqrteLUT[3109] = 16'hcc40;
RsqrteLUT[3110] = 16'hcc3d;
RsqrteLUT[3111] = 16'hcc3a;
RsqrteLUT[3112] = 16'hcc38;
RsqrteLUT[3113] = 16'hcc35;
RsqrteLUT[3114] = 16'hcc32;
RsqrteLUT[3115] = 16'hcc2f;
RsqrteLUT[3116] = 16'hcc2d;
RsqrteLUT[3117] = 16'hcc2a;
RsqrteLUT[3118] = 16'hcc28;
RsqrteLUT[3119] = 16'hcc25;
RsqrteLUT[3120] = 16'hcc23;
RsqrteLUT[3121] = 16'hcc20;
RsqrteLUT[3122] = 16'hcc1e;
RsqrteLUT[3123] = 16'hcc1c;
RsqrteLUT[3124] = 16'hcc19;
RsqrteLUT[3125] = 16'hcc17;
RsqrteLUT[3126] = 16'hcc15;
RsqrteLUT[3127] = 16'hcc13;
RsqrteLUT[3128] = 16'hcc10;
RsqrteLUT[3129] = 16'hcc0e;
RsqrteLUT[3130] = 16'hcc0c;
RsqrteLUT[3131] = 16'hcc0a;
RsqrteLUT[3132] = 16'hcc08;
RsqrteLUT[3133] = 16'hcc06;
RsqrteLUT[3134] = 16'hcc04;
RsqrteLUT[3135] = 16'hcc02;
RsqrteLUT[3136] = 16'hcc00;
RsqrteLUT[3137] = 16'hcbf8;
RsqrteLUT[3138] = 16'hcbf0;
RsqrteLUT[3139] = 16'hcbe8;
RsqrteLUT[3140] = 16'hcbe1;
RsqrteLUT[3141] = 16'hcbda;
RsqrteLUT[3142] = 16'hcbd3;
RsqrteLUT[3143] = 16'hcbcc;
RsqrteLUT[3144] = 16'hcbc5;
RsqrteLUT[3145] = 16'hcbbe;
RsqrteLUT[3146] = 16'hcbb8;
RsqrteLUT[3147] = 16'hcbb1;
RsqrteLUT[3148] = 16'hcbab;
RsqrteLUT[3149] = 16'hcba5;
RsqrteLUT[3150] = 16'hcb9f;
RsqrteLUT[3151] = 16'hcb99;
RsqrteLUT[3152] = 16'hcb93;
RsqrteLUT[3153] = 16'hcb8e;
RsqrteLUT[3154] = 16'hcb88;
RsqrteLUT[3155] = 16'hcb83;
RsqrteLUT[3156] = 16'hcb7d;
RsqrteLUT[3157] = 16'hcb78;
RsqrteLUT[3158] = 16'hcb73;
RsqrteLUT[3159] = 16'hcb6e;
RsqrteLUT[3160] = 16'hcb69;
RsqrteLUT[3161] = 16'hcb64;
RsqrteLUT[3162] = 16'hcb5f;
RsqrteLUT[3163] = 16'hcb5a;
RsqrteLUT[3164] = 16'hcb56;
RsqrteLUT[3165] = 16'hcb51;
RsqrteLUT[3166] = 16'hcb4c;
RsqrteLUT[3167] = 16'hcb48;
RsqrteLUT[3168] = 16'hcb44;
RsqrteLUT[3169] = 16'hcb3f;
RsqrteLUT[3170] = 16'hcb3b;
RsqrteLUT[3171] = 16'hcb37;
RsqrteLUT[3172] = 16'hcb33;
RsqrteLUT[3173] = 16'hcb2f;
RsqrteLUT[3174] = 16'hcb2b;
RsqrteLUT[3175] = 16'hcb27;
RsqrteLUT[3176] = 16'hcb23;
RsqrteLUT[3177] = 16'hcb1f;
RsqrteLUT[3178] = 16'hcb1b;
RsqrteLUT[3179] = 16'hcb17;
RsqrteLUT[3180] = 16'hcb14;
RsqrteLUT[3181] = 16'hcb10;
RsqrteLUT[3182] = 16'hcb0d;
RsqrteLUT[3183] = 16'hcb09;
RsqrteLUT[3184] = 16'hcb06;
RsqrteLUT[3185] = 16'hcb02;
RsqrteLUT[3186] = 16'hcaff;
RsqrteLUT[3187] = 16'hcafb;
RsqrteLUT[3188] = 16'hcaf8;
RsqrteLUT[3189] = 16'hcaf5;
RsqrteLUT[3190] = 16'hcaf2;
RsqrteLUT[3191] = 16'hcaee;
RsqrteLUT[3192] = 16'hcaeb;
RsqrteLUT[3193] = 16'hcae8;
RsqrteLUT[3194] = 16'hcae5;
RsqrteLUT[3195] = 16'hcae2;
RsqrteLUT[3196] = 16'hcadf;
RsqrteLUT[3197] = 16'hcadc;
RsqrteLUT[3198] = 16'hcad9;
RsqrteLUT[3199] = 16'hcad6;
RsqrteLUT[3200] = 16'hcad4;
RsqrteLUT[3201] = 16'hcace;
RsqrteLUT[3202] = 16'hcac9;
RsqrteLUT[3203] = 16'hcac3;
RsqrteLUT[3204] = 16'hcabe;
RsqrteLUT[3205] = 16'hcab9;
RsqrteLUT[3206] = 16'hcab4;
RsqrteLUT[3207] = 16'hcaaf;
RsqrteLUT[3208] = 16'hcaaa;
RsqrteLUT[3209] = 16'hcaa5;
RsqrteLUT[3210] = 16'hcaa1;
RsqrteLUT[3211] = 16'hca9c;
RsqrteLUT[3212] = 16'hca98;
RsqrteLUT[3213] = 16'hca94;
RsqrteLUT[3214] = 16'hca8f;
RsqrteLUT[3215] = 16'hca8b;
RsqrteLUT[3216] = 16'hca87;
RsqrteLUT[3217] = 16'hca83;
RsqrteLUT[3218] = 16'hca7f;
RsqrteLUT[3219] = 16'hca7b;
RsqrteLUT[3220] = 16'hca78;
RsqrteLUT[3221] = 16'hca74;
RsqrteLUT[3222] = 16'hca70;
RsqrteLUT[3223] = 16'hca6d;
RsqrteLUT[3224] = 16'hca69;
RsqrteLUT[3225] = 16'hca66;
RsqrteLUT[3226] = 16'hca62;
RsqrteLUT[3227] = 16'hca5f;
RsqrteLUT[3228] = 16'hca5b;
RsqrteLUT[3229] = 16'hca58;
RsqrteLUT[3230] = 16'hca55;
RsqrteLUT[3231] = 16'hca52;
RsqrteLUT[3232] = 16'hca4f;
RsqrteLUT[3233] = 16'hca4c;
RsqrteLUT[3234] = 16'hca49;
RsqrteLUT[3235] = 16'hca46;
RsqrteLUT[3236] = 16'hca43;
RsqrteLUT[3237] = 16'hca40;
RsqrteLUT[3238] = 16'hca3d;
RsqrteLUT[3239] = 16'hca3a;
RsqrteLUT[3240] = 16'hca38;
RsqrteLUT[3241] = 16'hca35;
RsqrteLUT[3242] = 16'hca32;
RsqrteLUT[3243] = 16'hca2f;
RsqrteLUT[3244] = 16'hca2d;
RsqrteLUT[3245] = 16'hca2a;
RsqrteLUT[3246] = 16'hca28;
RsqrteLUT[3247] = 16'hca25;
RsqrteLUT[3248] = 16'hca23;
RsqrteLUT[3249] = 16'hca20;
RsqrteLUT[3250] = 16'hca1e;
RsqrteLUT[3251] = 16'hca1c;
RsqrteLUT[3252] = 16'hca19;
RsqrteLUT[3253] = 16'hca17;
RsqrteLUT[3254] = 16'hca15;
RsqrteLUT[3255] = 16'hca13;
RsqrteLUT[3256] = 16'hca10;
RsqrteLUT[3257] = 16'hca0e;
RsqrteLUT[3258] = 16'hca0c;
RsqrteLUT[3259] = 16'hca0a;
RsqrteLUT[3260] = 16'hca08;
RsqrteLUT[3261] = 16'hca06;
RsqrteLUT[3262] = 16'hca04;
RsqrteLUT[3263] = 16'hca02;
RsqrteLUT[3264] = 16'hca00;
RsqrteLUT[3265] = 16'hc9f8;
RsqrteLUT[3266] = 16'hc9f0;
RsqrteLUT[3267] = 16'hc9e8;
RsqrteLUT[3268] = 16'hc9e1;
RsqrteLUT[3269] = 16'hc9da;
RsqrteLUT[3270] = 16'hc9d3;
RsqrteLUT[3271] = 16'hc9cc;
RsqrteLUT[3272] = 16'hc9c5;
RsqrteLUT[3273] = 16'hc9be;
RsqrteLUT[3274] = 16'hc9b8;
RsqrteLUT[3275] = 16'hc9b1;
RsqrteLUT[3276] = 16'hc9ab;
RsqrteLUT[3277] = 16'hc9a5;
RsqrteLUT[3278] = 16'hc99f;
RsqrteLUT[3279] = 16'hc999;
RsqrteLUT[3280] = 16'hc993;
RsqrteLUT[3281] = 16'hc98e;
RsqrteLUT[3282] = 16'hc988;
RsqrteLUT[3283] = 16'hc983;
RsqrteLUT[3284] = 16'hc97d;
RsqrteLUT[3285] = 16'hc978;
RsqrteLUT[3286] = 16'hc973;
RsqrteLUT[3287] = 16'hc96e;
RsqrteLUT[3288] = 16'hc969;
RsqrteLUT[3289] = 16'hc964;
RsqrteLUT[3290] = 16'hc95f;
RsqrteLUT[3291] = 16'hc95a;
RsqrteLUT[3292] = 16'hc956;
RsqrteLUT[3293] = 16'hc951;
RsqrteLUT[3294] = 16'hc94c;
RsqrteLUT[3295] = 16'hc948;
RsqrteLUT[3296] = 16'hc944;
RsqrteLUT[3297] = 16'hc93f;
RsqrteLUT[3298] = 16'hc93b;
RsqrteLUT[3299] = 16'hc937;
RsqrteLUT[3300] = 16'hc933;
RsqrteLUT[3301] = 16'hc92f;
RsqrteLUT[3302] = 16'hc92b;
RsqrteLUT[3303] = 16'hc927;
RsqrteLUT[3304] = 16'hc923;
RsqrteLUT[3305] = 16'hc91f;
RsqrteLUT[3306] = 16'hc91b;
RsqrteLUT[3307] = 16'hc917;
RsqrteLUT[3308] = 16'hc914;
RsqrteLUT[3309] = 16'hc910;
RsqrteLUT[3310] = 16'hc90d;
RsqrteLUT[3311] = 16'hc909;
RsqrteLUT[3312] = 16'hc906;
RsqrteLUT[3313] = 16'hc902;
RsqrteLUT[3314] = 16'hc8ff;
RsqrteLUT[3315] = 16'hc8fb;
RsqrteLUT[3316] = 16'hc8f8;
RsqrteLUT[3317] = 16'hc8f5;
RsqrteLUT[3318] = 16'hc8f2;
RsqrteLUT[3319] = 16'hc8ee;
RsqrteLUT[3320] = 16'hc8eb;
RsqrteLUT[3321] = 16'hc8e8;
RsqrteLUT[3322] = 16'hc8e5;
RsqrteLUT[3323] = 16'hc8e2;
RsqrteLUT[3324] = 16'hc8df;
RsqrteLUT[3325] = 16'hc8dc;
RsqrteLUT[3326] = 16'hc8d9;
RsqrteLUT[3327] = 16'hc8d6;
RsqrteLUT[3328] = 16'hc8d4;
RsqrteLUT[3329] = 16'hc8ce;
RsqrteLUT[3330] = 16'hc8c9;
RsqrteLUT[3331] = 16'hc8c3;
RsqrteLUT[3332] = 16'hc8be;
RsqrteLUT[3333] = 16'hc8b9;
RsqrteLUT[3334] = 16'hc8b4;
RsqrteLUT[3335] = 16'hc8af;
RsqrteLUT[3336] = 16'hc8aa;
RsqrteLUT[3337] = 16'hc8a5;
RsqrteLUT[3338] = 16'hc8a1;
RsqrteLUT[3339] = 16'hc89c;
RsqrteLUT[3340] = 16'hc898;
RsqrteLUT[3341] = 16'hc894;
RsqrteLUT[3342] = 16'hc88f;
RsqrteLUT[3343] = 16'hc88b;
RsqrteLUT[3344] = 16'hc887;
RsqrteLUT[3345] = 16'hc883;
RsqrteLUT[3346] = 16'hc87f;
RsqrteLUT[3347] = 16'hc87b;
RsqrteLUT[3348] = 16'hc878;
RsqrteLUT[3349] = 16'hc874;
RsqrteLUT[3350] = 16'hc870;
RsqrteLUT[3351] = 16'hc86d;
RsqrteLUT[3352] = 16'hc869;
RsqrteLUT[3353] = 16'hc866;
RsqrteLUT[3354] = 16'hc862;
RsqrteLUT[3355] = 16'hc85f;
RsqrteLUT[3356] = 16'hc85b;
RsqrteLUT[3357] = 16'hc858;
RsqrteLUT[3358] = 16'hc855;
RsqrteLUT[3359] = 16'hc852;
RsqrteLUT[3360] = 16'hc84f;
RsqrteLUT[3361] = 16'hc84c;
RsqrteLUT[3362] = 16'hc849;
RsqrteLUT[3363] = 16'hc846;
RsqrteLUT[3364] = 16'hc843;
RsqrteLUT[3365] = 16'hc840;
RsqrteLUT[3366] = 16'hc83d;
RsqrteLUT[3367] = 16'hc83a;
RsqrteLUT[3368] = 16'hc838;
RsqrteLUT[3369] = 16'hc835;
RsqrteLUT[3370] = 16'hc832;
RsqrteLUT[3371] = 16'hc82f;
RsqrteLUT[3372] = 16'hc82d;
RsqrteLUT[3373] = 16'hc82a;
RsqrteLUT[3374] = 16'hc828;
RsqrteLUT[3375] = 16'hc825;
RsqrteLUT[3376] = 16'hc823;
RsqrteLUT[3377] = 16'hc820;
RsqrteLUT[3378] = 16'hc81e;
RsqrteLUT[3379] = 16'hc81c;
RsqrteLUT[3380] = 16'hc819;
RsqrteLUT[3381] = 16'hc817;
RsqrteLUT[3382] = 16'hc815;
RsqrteLUT[3383] = 16'hc813;
RsqrteLUT[3384] = 16'hc810;
RsqrteLUT[3385] = 16'hc80e;
RsqrteLUT[3386] = 16'hc80c;
RsqrteLUT[3387] = 16'hc80a;
RsqrteLUT[3388] = 16'hc808;
RsqrteLUT[3389] = 16'hc806;
RsqrteLUT[3390] = 16'hc804;
RsqrteLUT[3391] = 16'hc802;
RsqrteLUT[3392] = 16'hc800;
RsqrteLUT[3393] = 16'hc7f8;
RsqrteLUT[3394] = 16'hc7f0;
RsqrteLUT[3395] = 16'hc7e8;
RsqrteLUT[3396] = 16'hc7e1;
RsqrteLUT[3397] = 16'hc7da;
RsqrteLUT[3398] = 16'hc7d3;
RsqrteLUT[3399] = 16'hc7cc;
RsqrteLUT[3400] = 16'hc7c5;
RsqrteLUT[3401] = 16'hc7be;
RsqrteLUT[3402] = 16'hc7b8;
RsqrteLUT[3403] = 16'hc7b1;
RsqrteLUT[3404] = 16'hc7ab;
RsqrteLUT[3405] = 16'hc7a5;
RsqrteLUT[3406] = 16'hc79f;
RsqrteLUT[3407] = 16'hc799;
RsqrteLUT[3408] = 16'hc793;
RsqrteLUT[3409] = 16'hc78e;
RsqrteLUT[3410] = 16'hc788;
RsqrteLUT[3411] = 16'hc783;
RsqrteLUT[3412] = 16'hc77d;
RsqrteLUT[3413] = 16'hc778;
RsqrteLUT[3414] = 16'hc773;
RsqrteLUT[3415] = 16'hc76e;
RsqrteLUT[3416] = 16'hc769;
RsqrteLUT[3417] = 16'hc764;
RsqrteLUT[3418] = 16'hc75f;
RsqrteLUT[3419] = 16'hc75a;
RsqrteLUT[3420] = 16'hc756;
RsqrteLUT[3421] = 16'hc751;
RsqrteLUT[3422] = 16'hc74c;
RsqrteLUT[3423] = 16'hc748;
RsqrteLUT[3424] = 16'hc744;
RsqrteLUT[3425] = 16'hc73f;
RsqrteLUT[3426] = 16'hc73b;
RsqrteLUT[3427] = 16'hc737;
RsqrteLUT[3428] = 16'hc733;
RsqrteLUT[3429] = 16'hc72f;
RsqrteLUT[3430] = 16'hc72b;
RsqrteLUT[3431] = 16'hc727;
RsqrteLUT[3432] = 16'hc723;
RsqrteLUT[3433] = 16'hc71f;
RsqrteLUT[3434] = 16'hc71b;
RsqrteLUT[3435] = 16'hc717;
RsqrteLUT[3436] = 16'hc714;
RsqrteLUT[3437] = 16'hc710;
RsqrteLUT[3438] = 16'hc70d;
RsqrteLUT[3439] = 16'hc709;
RsqrteLUT[3440] = 16'hc706;
RsqrteLUT[3441] = 16'hc702;
RsqrteLUT[3442] = 16'hc6ff;
RsqrteLUT[3443] = 16'hc6fb;
RsqrteLUT[3444] = 16'hc6f8;
RsqrteLUT[3445] = 16'hc6f5;
RsqrteLUT[3446] = 16'hc6f2;
RsqrteLUT[3447] = 16'hc6ee;
RsqrteLUT[3448] = 16'hc6eb;
RsqrteLUT[3449] = 16'hc6e8;
RsqrteLUT[3450] = 16'hc6e5;
RsqrteLUT[3451] = 16'hc6e2;
RsqrteLUT[3452] = 16'hc6df;
RsqrteLUT[3453] = 16'hc6dc;
RsqrteLUT[3454] = 16'hc6d9;
RsqrteLUT[3455] = 16'hc6d6;
RsqrteLUT[3456] = 16'hc6d4;
RsqrteLUT[3457] = 16'hc6ce;
RsqrteLUT[3458] = 16'hc6c9;
RsqrteLUT[3459] = 16'hc6c3;
RsqrteLUT[3460] = 16'hc6be;
RsqrteLUT[3461] = 16'hc6b9;
RsqrteLUT[3462] = 16'hc6b4;
RsqrteLUT[3463] = 16'hc6af;
RsqrteLUT[3464] = 16'hc6aa;
RsqrteLUT[3465] = 16'hc6a5;
RsqrteLUT[3466] = 16'hc6a1;
RsqrteLUT[3467] = 16'hc69c;
RsqrteLUT[3468] = 16'hc698;
RsqrteLUT[3469] = 16'hc694;
RsqrteLUT[3470] = 16'hc68f;
RsqrteLUT[3471] = 16'hc68b;
RsqrteLUT[3472] = 16'hc687;
RsqrteLUT[3473] = 16'hc683;
RsqrteLUT[3474] = 16'hc67f;
RsqrteLUT[3475] = 16'hc67b;
RsqrteLUT[3476] = 16'hc678;
RsqrteLUT[3477] = 16'hc674;
RsqrteLUT[3478] = 16'hc670;
RsqrteLUT[3479] = 16'hc66d;
RsqrteLUT[3480] = 16'hc669;
RsqrteLUT[3481] = 16'hc666;
RsqrteLUT[3482] = 16'hc662;
RsqrteLUT[3483] = 16'hc65f;
RsqrteLUT[3484] = 16'hc65b;
RsqrteLUT[3485] = 16'hc658;
RsqrteLUT[3486] = 16'hc655;
RsqrteLUT[3487] = 16'hc652;
RsqrteLUT[3488] = 16'hc64f;
RsqrteLUT[3489] = 16'hc64c;
RsqrteLUT[3490] = 16'hc649;
RsqrteLUT[3491] = 16'hc646;
RsqrteLUT[3492] = 16'hc643;
RsqrteLUT[3493] = 16'hc640;
RsqrteLUT[3494] = 16'hc63d;
RsqrteLUT[3495] = 16'hc63a;
RsqrteLUT[3496] = 16'hc638;
RsqrteLUT[3497] = 16'hc635;
RsqrteLUT[3498] = 16'hc632;
RsqrteLUT[3499] = 16'hc62f;
RsqrteLUT[3500] = 16'hc62d;
RsqrteLUT[3501] = 16'hc62a;
RsqrteLUT[3502] = 16'hc628;
RsqrteLUT[3503] = 16'hc625;
RsqrteLUT[3504] = 16'hc623;
RsqrteLUT[3505] = 16'hc620;
RsqrteLUT[3506] = 16'hc61e;
RsqrteLUT[3507] = 16'hc61c;
RsqrteLUT[3508] = 16'hc619;
RsqrteLUT[3509] = 16'hc617;
RsqrteLUT[3510] = 16'hc615;
RsqrteLUT[3511] = 16'hc613;
RsqrteLUT[3512] = 16'hc610;
RsqrteLUT[3513] = 16'hc60e;
RsqrteLUT[3514] = 16'hc60c;
RsqrteLUT[3515] = 16'hc60a;
RsqrteLUT[3516] = 16'hc608;
RsqrteLUT[3517] = 16'hc606;
RsqrteLUT[3518] = 16'hc604;
RsqrteLUT[3519] = 16'hc602;
RsqrteLUT[3520] = 16'hc600;
RsqrteLUT[3521] = 16'hc5f8;
RsqrteLUT[3522] = 16'hc5f0;
RsqrteLUT[3523] = 16'hc5e8;
RsqrteLUT[3524] = 16'hc5e1;
RsqrteLUT[3525] = 16'hc5da;
RsqrteLUT[3526] = 16'hc5d3;
RsqrteLUT[3527] = 16'hc5cc;
RsqrteLUT[3528] = 16'hc5c5;
RsqrteLUT[3529] = 16'hc5be;
RsqrteLUT[3530] = 16'hc5b8;
RsqrteLUT[3531] = 16'hc5b1;
RsqrteLUT[3532] = 16'hc5ab;
RsqrteLUT[3533] = 16'hc5a5;
RsqrteLUT[3534] = 16'hc59f;
RsqrteLUT[3535] = 16'hc599;
RsqrteLUT[3536] = 16'hc593;
RsqrteLUT[3537] = 16'hc58e;
RsqrteLUT[3538] = 16'hc588;
RsqrteLUT[3539] = 16'hc583;
RsqrteLUT[3540] = 16'hc57d;
RsqrteLUT[3541] = 16'hc578;
RsqrteLUT[3542] = 16'hc573;
RsqrteLUT[3543] = 16'hc56e;
RsqrteLUT[3544] = 16'hc569;
RsqrteLUT[3545] = 16'hc564;
RsqrteLUT[3546] = 16'hc55f;
RsqrteLUT[3547] = 16'hc55a;
RsqrteLUT[3548] = 16'hc556;
RsqrteLUT[3549] = 16'hc551;
RsqrteLUT[3550] = 16'hc54c;
RsqrteLUT[3551] = 16'hc548;
RsqrteLUT[3552] = 16'hc544;
RsqrteLUT[3553] = 16'hc53f;
RsqrteLUT[3554] = 16'hc53b;
RsqrteLUT[3555] = 16'hc537;
RsqrteLUT[3556] = 16'hc533;
RsqrteLUT[3557] = 16'hc52f;
RsqrteLUT[3558] = 16'hc52b;
RsqrteLUT[3559] = 16'hc527;
RsqrteLUT[3560] = 16'hc523;
RsqrteLUT[3561] = 16'hc51f;
RsqrteLUT[3562] = 16'hc51b;
RsqrteLUT[3563] = 16'hc517;
RsqrteLUT[3564] = 16'hc514;
RsqrteLUT[3565] = 16'hc510;
RsqrteLUT[3566] = 16'hc50d;
RsqrteLUT[3567] = 16'hc509;
RsqrteLUT[3568] = 16'hc506;
RsqrteLUT[3569] = 16'hc502;
RsqrteLUT[3570] = 16'hc4ff;
RsqrteLUT[3571] = 16'hc4fb;
RsqrteLUT[3572] = 16'hc4f8;
RsqrteLUT[3573] = 16'hc4f5;
RsqrteLUT[3574] = 16'hc4f2;
RsqrteLUT[3575] = 16'hc4ee;
RsqrteLUT[3576] = 16'hc4eb;
RsqrteLUT[3577] = 16'hc4e8;
RsqrteLUT[3578] = 16'hc4e5;
RsqrteLUT[3579] = 16'hc4e2;
RsqrteLUT[3580] = 16'hc4df;
RsqrteLUT[3581] = 16'hc4dc;
RsqrteLUT[3582] = 16'hc4d9;
RsqrteLUT[3583] = 16'hc4d6;
RsqrteLUT[3584] = 16'hc4d4;
RsqrteLUT[3585] = 16'hc4ce;
RsqrteLUT[3586] = 16'hc4c9;
RsqrteLUT[3587] = 16'hc4c3;
RsqrteLUT[3588] = 16'hc4be;
RsqrteLUT[3589] = 16'hc4b9;
RsqrteLUT[3590] = 16'hc4b4;
RsqrteLUT[3591] = 16'hc4af;
RsqrteLUT[3592] = 16'hc4aa;
RsqrteLUT[3593] = 16'hc4a5;
RsqrteLUT[3594] = 16'hc4a1;
RsqrteLUT[3595] = 16'hc49c;
RsqrteLUT[3596] = 16'hc498;
RsqrteLUT[3597] = 16'hc494;
RsqrteLUT[3598] = 16'hc48f;
RsqrteLUT[3599] = 16'hc48b;
RsqrteLUT[3600] = 16'hc487;
RsqrteLUT[3601] = 16'hc483;
RsqrteLUT[3602] = 16'hc47f;
RsqrteLUT[3603] = 16'hc47b;
RsqrteLUT[3604] = 16'hc478;
RsqrteLUT[3605] = 16'hc474;
RsqrteLUT[3606] = 16'hc470;
RsqrteLUT[3607] = 16'hc46d;
RsqrteLUT[3608] = 16'hc469;
RsqrteLUT[3609] = 16'hc466;
RsqrteLUT[3610] = 16'hc462;
RsqrteLUT[3611] = 16'hc45f;
RsqrteLUT[3612] = 16'hc45b;
RsqrteLUT[3613] = 16'hc458;
RsqrteLUT[3614] = 16'hc455;
RsqrteLUT[3615] = 16'hc452;
RsqrteLUT[3616] = 16'hc44f;
RsqrteLUT[3617] = 16'hc44c;
RsqrteLUT[3618] = 16'hc449;
RsqrteLUT[3619] = 16'hc446;
RsqrteLUT[3620] = 16'hc443;
RsqrteLUT[3621] = 16'hc440;
RsqrteLUT[3622] = 16'hc43d;
RsqrteLUT[3623] = 16'hc43a;
RsqrteLUT[3624] = 16'hc438;
RsqrteLUT[3625] = 16'hc435;
RsqrteLUT[3626] = 16'hc432;
RsqrteLUT[3627] = 16'hc42f;
RsqrteLUT[3628] = 16'hc42d;
RsqrteLUT[3629] = 16'hc42a;
RsqrteLUT[3630] = 16'hc428;
RsqrteLUT[3631] = 16'hc425;
RsqrteLUT[3632] = 16'hc423;
RsqrteLUT[3633] = 16'hc420;
RsqrteLUT[3634] = 16'hc41e;
RsqrteLUT[3635] = 16'hc41c;
RsqrteLUT[3636] = 16'hc419;
RsqrteLUT[3637] = 16'hc417;
RsqrteLUT[3638] = 16'hc415;
RsqrteLUT[3639] = 16'hc413;
RsqrteLUT[3640] = 16'hc410;
RsqrteLUT[3641] = 16'hc40e;
RsqrteLUT[3642] = 16'hc40c;
RsqrteLUT[3643] = 16'hc40a;
RsqrteLUT[3644] = 16'hc408;
RsqrteLUT[3645] = 16'hc406;
RsqrteLUT[3646] = 16'hc404;
RsqrteLUT[3647] = 16'hc402;
RsqrteLUT[3648] = 16'hc400;
RsqrteLUT[3649] = 16'hc3f8;
RsqrteLUT[3650] = 16'hc3f0;
RsqrteLUT[3651] = 16'hc3e8;
RsqrteLUT[3652] = 16'hc3e1;
RsqrteLUT[3653] = 16'hc3da;
RsqrteLUT[3654] = 16'hc3d3;
RsqrteLUT[3655] = 16'hc3cc;
RsqrteLUT[3656] = 16'hc3c5;
RsqrteLUT[3657] = 16'hc3be;
RsqrteLUT[3658] = 16'hc3b8;
RsqrteLUT[3659] = 16'hc3b1;
RsqrteLUT[3660] = 16'hc3ab;
RsqrteLUT[3661] = 16'hc3a5;
RsqrteLUT[3662] = 16'hc39f;
RsqrteLUT[3663] = 16'hc399;
RsqrteLUT[3664] = 16'hc393;
RsqrteLUT[3665] = 16'hc38e;
RsqrteLUT[3666] = 16'hc388;
RsqrteLUT[3667] = 16'hc383;
RsqrteLUT[3668] = 16'hc37d;
RsqrteLUT[3669] = 16'hc378;
RsqrteLUT[3670] = 16'hc373;
RsqrteLUT[3671] = 16'hc36e;
RsqrteLUT[3672] = 16'hc369;
RsqrteLUT[3673] = 16'hc364;
RsqrteLUT[3674] = 16'hc35f;
RsqrteLUT[3675] = 16'hc35a;
RsqrteLUT[3676] = 16'hc356;
RsqrteLUT[3677] = 16'hc351;
RsqrteLUT[3678] = 16'hc34c;
RsqrteLUT[3679] = 16'hc348;
RsqrteLUT[3680] = 16'hc344;
RsqrteLUT[3681] = 16'hc33f;
RsqrteLUT[3682] = 16'hc33b;
RsqrteLUT[3683] = 16'hc337;
RsqrteLUT[3684] = 16'hc333;
RsqrteLUT[3685] = 16'hc32f;
RsqrteLUT[3686] = 16'hc32b;
RsqrteLUT[3687] = 16'hc327;
RsqrteLUT[3688] = 16'hc323;
RsqrteLUT[3689] = 16'hc31f;
RsqrteLUT[3690] = 16'hc31b;
RsqrteLUT[3691] = 16'hc317;
RsqrteLUT[3692] = 16'hc314;
RsqrteLUT[3693] = 16'hc310;
RsqrteLUT[3694] = 16'hc30d;
RsqrteLUT[3695] = 16'hc309;
RsqrteLUT[3696] = 16'hc306;
RsqrteLUT[3697] = 16'hc302;
RsqrteLUT[3698] = 16'hc2ff;
RsqrteLUT[3699] = 16'hc2fb;
RsqrteLUT[3700] = 16'hc2f8;
RsqrteLUT[3701] = 16'hc2f5;
RsqrteLUT[3702] = 16'hc2f2;
RsqrteLUT[3703] = 16'hc2ee;
RsqrteLUT[3704] = 16'hc2eb;
RsqrteLUT[3705] = 16'hc2e8;
RsqrteLUT[3706] = 16'hc2e5;
RsqrteLUT[3707] = 16'hc2e2;
RsqrteLUT[3708] = 16'hc2df;
RsqrteLUT[3709] = 16'hc2dc;
RsqrteLUT[3710] = 16'hc2d9;
RsqrteLUT[3711] = 16'hc2d6;
RsqrteLUT[3712] = 16'hc2d4;
RsqrteLUT[3713] = 16'hc2ce;
RsqrteLUT[3714] = 16'hc2c9;
RsqrteLUT[3715] = 16'hc2c3;
RsqrteLUT[3716] = 16'hc2be;
RsqrteLUT[3717] = 16'hc2b9;
RsqrteLUT[3718] = 16'hc2b4;
RsqrteLUT[3719] = 16'hc2af;
RsqrteLUT[3720] = 16'hc2aa;
RsqrteLUT[3721] = 16'hc2a5;
RsqrteLUT[3722] = 16'hc2a1;
RsqrteLUT[3723] = 16'hc29c;
RsqrteLUT[3724] = 16'hc298;
RsqrteLUT[3725] = 16'hc294;
RsqrteLUT[3726] = 16'hc28f;
RsqrteLUT[3727] = 16'hc28b;
RsqrteLUT[3728] = 16'hc287;
RsqrteLUT[3729] = 16'hc283;
RsqrteLUT[3730] = 16'hc27f;
RsqrteLUT[3731] = 16'hc27b;
RsqrteLUT[3732] = 16'hc278;
RsqrteLUT[3733] = 16'hc274;
RsqrteLUT[3734] = 16'hc270;
RsqrteLUT[3735] = 16'hc26d;
RsqrteLUT[3736] = 16'hc269;
RsqrteLUT[3737] = 16'hc266;
RsqrteLUT[3738] = 16'hc262;
RsqrteLUT[3739] = 16'hc25f;
RsqrteLUT[3740] = 16'hc25b;
RsqrteLUT[3741] = 16'hc258;
RsqrteLUT[3742] = 16'hc255;
RsqrteLUT[3743] = 16'hc252;
RsqrteLUT[3744] = 16'hc24f;
RsqrteLUT[3745] = 16'hc24c;
RsqrteLUT[3746] = 16'hc249;
RsqrteLUT[3747] = 16'hc246;
RsqrteLUT[3748] = 16'hc243;
RsqrteLUT[3749] = 16'hc240;
RsqrteLUT[3750] = 16'hc23d;
RsqrteLUT[3751] = 16'hc23a;
RsqrteLUT[3752] = 16'hc238;
RsqrteLUT[3753] = 16'hc235;
RsqrteLUT[3754] = 16'hc232;
RsqrteLUT[3755] = 16'hc22f;
RsqrteLUT[3756] = 16'hc22d;
RsqrteLUT[3757] = 16'hc22a;
RsqrteLUT[3758] = 16'hc228;
RsqrteLUT[3759] = 16'hc225;
RsqrteLUT[3760] = 16'hc223;
RsqrteLUT[3761] = 16'hc220;
RsqrteLUT[3762] = 16'hc21e;
RsqrteLUT[3763] = 16'hc21c;
RsqrteLUT[3764] = 16'hc219;
RsqrteLUT[3765] = 16'hc217;
RsqrteLUT[3766] = 16'hc215;
RsqrteLUT[3767] = 16'hc213;
RsqrteLUT[3768] = 16'hc210;
RsqrteLUT[3769] = 16'hc20e;
RsqrteLUT[3770] = 16'hc20c;
RsqrteLUT[3771] = 16'hc20a;
RsqrteLUT[3772] = 16'hc208;
RsqrteLUT[3773] = 16'hc206;
RsqrteLUT[3774] = 16'hc204;
RsqrteLUT[3775] = 16'hc202;
RsqrteLUT[3776] = 16'hc200;
RsqrteLUT[3777] = 16'hc1f8;
RsqrteLUT[3778] = 16'hc1f0;
RsqrteLUT[3779] = 16'hc1e8;
RsqrteLUT[3780] = 16'hc1e1;
RsqrteLUT[3781] = 16'hc1da;
RsqrteLUT[3782] = 16'hc1d3;
RsqrteLUT[3783] = 16'hc1cc;
RsqrteLUT[3784] = 16'hc1c5;
RsqrteLUT[3785] = 16'hc1be;
RsqrteLUT[3786] = 16'hc1b8;
RsqrteLUT[3787] = 16'hc1b1;
RsqrteLUT[3788] = 16'hc1ab;
RsqrteLUT[3789] = 16'hc1a5;
RsqrteLUT[3790] = 16'hc19f;
RsqrteLUT[3791] = 16'hc199;
RsqrteLUT[3792] = 16'hc193;
RsqrteLUT[3793] = 16'hc18e;
RsqrteLUT[3794] = 16'hc188;
RsqrteLUT[3795] = 16'hc183;
RsqrteLUT[3796] = 16'hc17d;
RsqrteLUT[3797] = 16'hc178;
RsqrteLUT[3798] = 16'hc173;
RsqrteLUT[3799] = 16'hc16e;
RsqrteLUT[3800] = 16'hc169;
RsqrteLUT[3801] = 16'hc164;
RsqrteLUT[3802] = 16'hc15f;
RsqrteLUT[3803] = 16'hc15a;
RsqrteLUT[3804] = 16'hc156;
RsqrteLUT[3805] = 16'hc151;
RsqrteLUT[3806] = 16'hc14c;
RsqrteLUT[3807] = 16'hc148;
RsqrteLUT[3808] = 16'hc144;
RsqrteLUT[3809] = 16'hc13f;
RsqrteLUT[3810] = 16'hc13b;
RsqrteLUT[3811] = 16'hc137;
RsqrteLUT[3812] = 16'hc133;
RsqrteLUT[3813] = 16'hc12f;
RsqrteLUT[3814] = 16'hc12b;
RsqrteLUT[3815] = 16'hc127;
RsqrteLUT[3816] = 16'hc123;
RsqrteLUT[3817] = 16'hc11f;
RsqrteLUT[3818] = 16'hc11b;
RsqrteLUT[3819] = 16'hc117;
RsqrteLUT[3820] = 16'hc114;
RsqrteLUT[3821] = 16'hc110;
RsqrteLUT[3822] = 16'hc10d;
RsqrteLUT[3823] = 16'hc109;
RsqrteLUT[3824] = 16'hc106;
RsqrteLUT[3825] = 16'hc102;
RsqrteLUT[3826] = 16'hc0ff;
RsqrteLUT[3827] = 16'hc0fb;
RsqrteLUT[3828] = 16'hc0f8;
RsqrteLUT[3829] = 16'hc0f5;
RsqrteLUT[3830] = 16'hc0f2;
RsqrteLUT[3831] = 16'hc0ee;
RsqrteLUT[3832] = 16'hc0eb;
RsqrteLUT[3833] = 16'hc0e8;
RsqrteLUT[3834] = 16'hc0e5;
RsqrteLUT[3835] = 16'hc0e2;
RsqrteLUT[3836] = 16'hc0df;
RsqrteLUT[3837] = 16'hc0dc;
RsqrteLUT[3838] = 16'hc0d9;
RsqrteLUT[3839] = 16'hc0d6;
RsqrteLUT[3840] = 16'hc0d4;
RsqrteLUT[3841] = 16'hc0ce;
RsqrteLUT[3842] = 16'hc0c9;
RsqrteLUT[3843] = 16'hc0c3;
RsqrteLUT[3844] = 16'hc0be;
RsqrteLUT[3845] = 16'hc0b9;
RsqrteLUT[3846] = 16'hc0b4;
RsqrteLUT[3847] = 16'hc0af;
RsqrteLUT[3848] = 16'hc0aa;
RsqrteLUT[3849] = 16'hc0a5;
RsqrteLUT[3850] = 16'hc0a1;
RsqrteLUT[3851] = 16'hc09c;
RsqrteLUT[3852] = 16'hc098;
RsqrteLUT[3853] = 16'hc094;
RsqrteLUT[3854] = 16'hc08f;
RsqrteLUT[3855] = 16'hc08b;
RsqrteLUT[3856] = 16'hc087;
RsqrteLUT[3857] = 16'hc083;
RsqrteLUT[3858] = 16'hc07f;
RsqrteLUT[3859] = 16'hc07b;
RsqrteLUT[3860] = 16'hc078;
RsqrteLUT[3861] = 16'hc074;
RsqrteLUT[3862] = 16'hc070;
RsqrteLUT[3863] = 16'hc06d;
RsqrteLUT[3864] = 16'hc069;
RsqrteLUT[3865] = 16'hc066;
RsqrteLUT[3866] = 16'hc062;
RsqrteLUT[3867] = 16'hc05f;
RsqrteLUT[3868] = 16'hc05b;
RsqrteLUT[3869] = 16'hc058;
RsqrteLUT[3870] = 16'hc055;
RsqrteLUT[3871] = 16'hc052;
RsqrteLUT[3872] = 16'hc04f;
RsqrteLUT[3873] = 16'hc04c;
RsqrteLUT[3874] = 16'hc049;
RsqrteLUT[3875] = 16'hc046;
RsqrteLUT[3876] = 16'hc043;
RsqrteLUT[3877] = 16'hc040;
RsqrteLUT[3878] = 16'hc03d;
RsqrteLUT[3879] = 16'hc03a;
RsqrteLUT[3880] = 16'hc038;
RsqrteLUT[3881] = 16'hc035;
RsqrteLUT[3882] = 16'hc032;
RsqrteLUT[3883] = 16'hc02f;
RsqrteLUT[3884] = 16'hc02d;
RsqrteLUT[3885] = 16'hc02a;
RsqrteLUT[3886] = 16'hc028;
RsqrteLUT[3887] = 16'hc025;
RsqrteLUT[3888] = 16'hc023;
RsqrteLUT[3889] = 16'hc020;
RsqrteLUT[3890] = 16'hc01e;
RsqrteLUT[3891] = 16'hc01c;
RsqrteLUT[3892] = 16'hc019;
RsqrteLUT[3893] = 16'hc017;
RsqrteLUT[3894] = 16'hc015;
RsqrteLUT[3895] = 16'hc013;
RsqrteLUT[3896] = 16'hc010;
RsqrteLUT[3897] = 16'hc00e;
RsqrteLUT[3898] = 16'hc00c;
RsqrteLUT[3899] = 16'hc00a;
RsqrteLUT[3900] = 16'hc008;
RsqrteLUT[3901] = 16'hc006;
RsqrteLUT[3902] = 16'hc004;
RsqrteLUT[3903] = 16'hc002;
RsqrteLUT[3904] = 16'hc000;
RsqrteLUT[3905] = 16'hbff8;
RsqrteLUT[3906] = 16'hbff0;
RsqrteLUT[3907] = 16'hbfe8;
RsqrteLUT[3908] = 16'hbfe1;
RsqrteLUT[3909] = 16'hbfda;
RsqrteLUT[3910] = 16'hbfd3;
RsqrteLUT[3911] = 16'hbfcc;
RsqrteLUT[3912] = 16'hbfc5;
RsqrteLUT[3913] = 16'hbfbe;
RsqrteLUT[3914] = 16'hbfb8;
RsqrteLUT[3915] = 16'hbfb1;
RsqrteLUT[3916] = 16'hbfab;
RsqrteLUT[3917] = 16'hbfa5;
RsqrteLUT[3918] = 16'hbf9f;
RsqrteLUT[3919] = 16'hbf99;
RsqrteLUT[3920] = 16'hbf93;
RsqrteLUT[3921] = 16'hbf8e;
RsqrteLUT[3922] = 16'hbf88;
RsqrteLUT[3923] = 16'hbf83;
RsqrteLUT[3924] = 16'hbf7d;
RsqrteLUT[3925] = 16'hbf78;
RsqrteLUT[3926] = 16'hbf73;
RsqrteLUT[3927] = 16'hbf6e;
RsqrteLUT[3928] = 16'hbf69;
RsqrteLUT[3929] = 16'hbf64;
RsqrteLUT[3930] = 16'hbf5f;
RsqrteLUT[3931] = 16'hbf5a;
RsqrteLUT[3932] = 16'hbf56;
RsqrteLUT[3933] = 16'hbf51;
RsqrteLUT[3934] = 16'hbf4c;
RsqrteLUT[3935] = 16'hbf48;
RsqrteLUT[3936] = 16'hbf44;
RsqrteLUT[3937] = 16'hbf3f;
RsqrteLUT[3938] = 16'hbf3b;
RsqrteLUT[3939] = 16'hbf37;
RsqrteLUT[3940] = 16'hbf33;
RsqrteLUT[3941] = 16'hbf2f;
RsqrteLUT[3942] = 16'hbf2b;
RsqrteLUT[3943] = 16'hbf27;
RsqrteLUT[3944] = 16'hbf23;
RsqrteLUT[3945] = 16'hbf1f;
RsqrteLUT[3946] = 16'hbf1b;
RsqrteLUT[3947] = 16'hbf17;
RsqrteLUT[3948] = 16'hbf14;
RsqrteLUT[3949] = 16'hbf10;
RsqrteLUT[3950] = 16'hbf0d;
RsqrteLUT[3951] = 16'hbf09;
RsqrteLUT[3952] = 16'hbf06;
RsqrteLUT[3953] = 16'hbf02;
RsqrteLUT[3954] = 16'hbeff;
RsqrteLUT[3955] = 16'hbefb;
RsqrteLUT[3956] = 16'hbef8;
RsqrteLUT[3957] = 16'hbef5;
RsqrteLUT[3958] = 16'hbef2;
RsqrteLUT[3959] = 16'hbeee;
RsqrteLUT[3960] = 16'hbeeb;
RsqrteLUT[3961] = 16'hbee8;
RsqrteLUT[3962] = 16'hbee5;
RsqrteLUT[3963] = 16'hbee2;
RsqrteLUT[3964] = 16'hbedf;
RsqrteLUT[3965] = 16'hbedc;
RsqrteLUT[3966] = 16'hbed9;
RsqrteLUT[3967] = 16'hbed6;
RsqrteLUT[3968] = 16'hbed4;
RsqrteLUT[3969] = 16'hbece;
RsqrteLUT[3970] = 16'hbec9;
RsqrteLUT[3971] = 16'hbec3;
RsqrteLUT[3972] = 16'hbebe;
RsqrteLUT[3973] = 16'hbeb9;
RsqrteLUT[3974] = 16'hbeb4;
RsqrteLUT[3975] = 16'hbeaf;
RsqrteLUT[3976] = 16'hbeaa;
RsqrteLUT[3977] = 16'hbea5;
RsqrteLUT[3978] = 16'hbea1;
RsqrteLUT[3979] = 16'hbe9c;
RsqrteLUT[3980] = 16'hbe98;
RsqrteLUT[3981] = 16'hbe94;
RsqrteLUT[3982] = 16'hbe8f;
RsqrteLUT[3983] = 16'hbe8b;
RsqrteLUT[3984] = 16'hbe87;
RsqrteLUT[3985] = 16'hbe83;
RsqrteLUT[3986] = 16'hbe7f;
RsqrteLUT[3987] = 16'hbe7b;
RsqrteLUT[3988] = 16'hbe78;
RsqrteLUT[3989] = 16'hbe74;
RsqrteLUT[3990] = 16'hbe70;
RsqrteLUT[3991] = 16'hbe6d;
RsqrteLUT[3992] = 16'hbe69;
RsqrteLUT[3993] = 16'hbe66;
RsqrteLUT[3994] = 16'hbe62;
RsqrteLUT[3995] = 16'hbe5f;
RsqrteLUT[3996] = 16'hbe5b;
RsqrteLUT[3997] = 16'hbe58;
RsqrteLUT[3998] = 16'hbe55;
RsqrteLUT[3999] = 16'hbe52;
RsqrteLUT[4000] = 16'hbe4f;
RsqrteLUT[4001] = 16'hbe4c;
RsqrteLUT[4002] = 16'hbe49;
RsqrteLUT[4003] = 16'hbe46;
RsqrteLUT[4004] = 16'hbe43;
RsqrteLUT[4005] = 16'hbe40;
RsqrteLUT[4006] = 16'hbe3d;
RsqrteLUT[4007] = 16'hbe3a;
RsqrteLUT[4008] = 16'hbe38;
RsqrteLUT[4009] = 16'hbe35;
RsqrteLUT[4010] = 16'hbe32;
RsqrteLUT[4011] = 16'hbe2f;
RsqrteLUT[4012] = 16'hbe2d;
RsqrteLUT[4013] = 16'hbe2a;
RsqrteLUT[4014] = 16'hbe28;
RsqrteLUT[4015] = 16'hbe25;
RsqrteLUT[4016] = 16'hbe23;
RsqrteLUT[4017] = 16'hbe20;
RsqrteLUT[4018] = 16'hbe1e;
RsqrteLUT[4019] = 16'hbe1c;
RsqrteLUT[4020] = 16'hbe19;
RsqrteLUT[4021] = 16'hbe17;
RsqrteLUT[4022] = 16'hbe15;
RsqrteLUT[4023] = 16'hbe13;
RsqrteLUT[4024] = 16'hbe10;
RsqrteLUT[4025] = 16'hbe0e;
RsqrteLUT[4026] = 16'hbe0c;
RsqrteLUT[4027] = 16'hbe0a;
RsqrteLUT[4028] = 16'hbe08;
RsqrteLUT[4029] = 16'hbe06;
RsqrteLUT[4030] = 16'hbe04;
RsqrteLUT[4031] = 16'hbe02;
RsqrteLUT[4032] = 16'hbe00;
RsqrteLUT[4033] = 16'hbdf8;
RsqrteLUT[4034] = 16'hbdf0;
RsqrteLUT[4035] = 16'hbde8;
RsqrteLUT[4036] = 16'hbde1;
RsqrteLUT[4037] = 16'hbdda;
RsqrteLUT[4038] = 16'hbdd3;
RsqrteLUT[4039] = 16'hbdcc;
RsqrteLUT[4040] = 16'hbdc5;
RsqrteLUT[4041] = 16'hbdbe;
RsqrteLUT[4042] = 16'hbdb8;
RsqrteLUT[4043] = 16'hbdb1;
RsqrteLUT[4044] = 16'hbdab;
RsqrteLUT[4045] = 16'hbda5;
RsqrteLUT[4046] = 16'hbd9f;
RsqrteLUT[4047] = 16'hbd99;
RsqrteLUT[4048] = 16'hbd93;
RsqrteLUT[4049] = 16'hbd8e;
RsqrteLUT[4050] = 16'hbd88;
RsqrteLUT[4051] = 16'hbd83;
RsqrteLUT[4052] = 16'hbd7d;
RsqrteLUT[4053] = 16'hbd78;
RsqrteLUT[4054] = 16'hbd73;
RsqrteLUT[4055] = 16'hbd6e;
RsqrteLUT[4056] = 16'hbd69;
RsqrteLUT[4057] = 16'hbd64;
RsqrteLUT[4058] = 16'hbd5f;
RsqrteLUT[4059] = 16'hbd5a;
RsqrteLUT[4060] = 16'hbd56;
RsqrteLUT[4061] = 16'hbd51;
RsqrteLUT[4062] = 16'hbd4c;
RsqrteLUT[4063] = 16'hbd48;
RsqrteLUT[4064] = 16'hbd44;
RsqrteLUT[4065] = 16'hbd3f;
RsqrteLUT[4066] = 16'hbd3b;
RsqrteLUT[4067] = 16'hbd37;
RsqrteLUT[4068] = 16'hbd33;
RsqrteLUT[4069] = 16'hbd2f;
RsqrteLUT[4070] = 16'hbd2b;
RsqrteLUT[4071] = 16'hbd27;
RsqrteLUT[4072] = 16'hbd23;
RsqrteLUT[4073] = 16'hbd1f;
RsqrteLUT[4074] = 16'hbd1b;
RsqrteLUT[4075] = 16'hbd17;
RsqrteLUT[4076] = 16'hbd14;
RsqrteLUT[4077] = 16'hbd10;
RsqrteLUT[4078] = 16'hbd0d;
RsqrteLUT[4079] = 16'hbd09;
RsqrteLUT[4080] = 16'hbd06;
RsqrteLUT[4081] = 16'hbd02;
RsqrteLUT[4082] = 16'hbcff;
RsqrteLUT[4083] = 16'hbcfb;
RsqrteLUT[4084] = 16'hbcf8;
RsqrteLUT[4085] = 16'hbcf5;
RsqrteLUT[4086] = 16'hbcf2;
RsqrteLUT[4087] = 16'hbcee;
RsqrteLUT[4088] = 16'hbceb;
RsqrteLUT[4089] = 16'hbce8;
RsqrteLUT[4090] = 16'hbce5;
RsqrteLUT[4091] = 16'hbce2;
RsqrteLUT[4092] = 16'hbcdf;
RsqrteLUT[4093] = 16'hbcdc;
RsqrteLUT[4094] = 16'hbcd9;
RsqrteLUT[4095] = 16'hbcd6;
RsqrteLUT[4096] = 16'hbcd4;
RsqrteLUT[4097] = 16'hbcce;
RsqrteLUT[4098] = 16'hbcc9;
RsqrteLUT[4099] = 16'hbcc3;
RsqrteLUT[4100] = 16'hbcbe;
RsqrteLUT[4101] = 16'hbcb9;
RsqrteLUT[4102] = 16'hbcb4;
RsqrteLUT[4103] = 16'hbcaf;
RsqrteLUT[4104] = 16'hbcaa;
RsqrteLUT[4105] = 16'hbca5;
RsqrteLUT[4106] = 16'hbca1;
RsqrteLUT[4107] = 16'hbc9c;
RsqrteLUT[4108] = 16'hbc98;
RsqrteLUT[4109] = 16'hbc94;
RsqrteLUT[4110] = 16'hbc8f;
RsqrteLUT[4111] = 16'hbc8b;
RsqrteLUT[4112] = 16'hbc87;
RsqrteLUT[4113] = 16'hbc83;
RsqrteLUT[4114] = 16'hbc7f;
RsqrteLUT[4115] = 16'hbc7b;
RsqrteLUT[4116] = 16'hbc78;
RsqrteLUT[4117] = 16'hbc74;
RsqrteLUT[4118] = 16'hbc70;
RsqrteLUT[4119] = 16'hbc6d;
RsqrteLUT[4120] = 16'hbc69;
RsqrteLUT[4121] = 16'hbc66;
RsqrteLUT[4122] = 16'hbc62;
RsqrteLUT[4123] = 16'hbc5f;
RsqrteLUT[4124] = 16'hbc5b;
RsqrteLUT[4125] = 16'hbc58;
RsqrteLUT[4126] = 16'hbc55;
RsqrteLUT[4127] = 16'hbc52;
RsqrteLUT[4128] = 16'hbc4f;
RsqrteLUT[4129] = 16'hbc4c;
RsqrteLUT[4130] = 16'hbc49;
RsqrteLUT[4131] = 16'hbc46;
RsqrteLUT[4132] = 16'hbc43;
RsqrteLUT[4133] = 16'hbc40;
RsqrteLUT[4134] = 16'hbc3d;
RsqrteLUT[4135] = 16'hbc3a;
RsqrteLUT[4136] = 16'hbc38;
RsqrteLUT[4137] = 16'hbc35;
RsqrteLUT[4138] = 16'hbc32;
RsqrteLUT[4139] = 16'hbc2f;
RsqrteLUT[4140] = 16'hbc2d;
RsqrteLUT[4141] = 16'hbc2a;
RsqrteLUT[4142] = 16'hbc28;
RsqrteLUT[4143] = 16'hbc25;
RsqrteLUT[4144] = 16'hbc23;
RsqrteLUT[4145] = 16'hbc20;
RsqrteLUT[4146] = 16'hbc1e;
RsqrteLUT[4147] = 16'hbc1c;
RsqrteLUT[4148] = 16'hbc19;
RsqrteLUT[4149] = 16'hbc17;
RsqrteLUT[4150] = 16'hbc15;
RsqrteLUT[4151] = 16'hbc13;
RsqrteLUT[4152] = 16'hbc10;
RsqrteLUT[4153] = 16'hbc0e;
RsqrteLUT[4154] = 16'hbc0c;
RsqrteLUT[4155] = 16'hbc0a;
RsqrteLUT[4156] = 16'hbc08;
RsqrteLUT[4157] = 16'hbc06;
RsqrteLUT[4158] = 16'hbc04;
RsqrteLUT[4159] = 16'hbc02;
RsqrteLUT[4160] = 16'hbc00;
RsqrteLUT[4161] = 16'hbbf8;
RsqrteLUT[4162] = 16'hbbf0;
RsqrteLUT[4163] = 16'hbbe8;
RsqrteLUT[4164] = 16'hbbe1;
RsqrteLUT[4165] = 16'hbbda;
RsqrteLUT[4166] = 16'hbbd3;
RsqrteLUT[4167] = 16'hbbcc;
RsqrteLUT[4168] = 16'hbbc5;
RsqrteLUT[4169] = 16'hbbbe;
RsqrteLUT[4170] = 16'hbbb8;
RsqrteLUT[4171] = 16'hbbb1;
RsqrteLUT[4172] = 16'hbbab;
RsqrteLUT[4173] = 16'hbba5;
RsqrteLUT[4174] = 16'hbb9f;
RsqrteLUT[4175] = 16'hbb99;
RsqrteLUT[4176] = 16'hbb93;
RsqrteLUT[4177] = 16'hbb8e;
RsqrteLUT[4178] = 16'hbb88;
RsqrteLUT[4179] = 16'hbb83;
RsqrteLUT[4180] = 16'hbb7d;
RsqrteLUT[4181] = 16'hbb78;
RsqrteLUT[4182] = 16'hbb73;
RsqrteLUT[4183] = 16'hbb6e;
RsqrteLUT[4184] = 16'hbb69;
RsqrteLUT[4185] = 16'hbb64;
RsqrteLUT[4186] = 16'hbb5f;
RsqrteLUT[4187] = 16'hbb5a;
RsqrteLUT[4188] = 16'hbb56;
RsqrteLUT[4189] = 16'hbb51;
RsqrteLUT[4190] = 16'hbb4c;
RsqrteLUT[4191] = 16'hbb48;
RsqrteLUT[4192] = 16'hbb44;
RsqrteLUT[4193] = 16'hbb3f;
RsqrteLUT[4194] = 16'hbb3b;
RsqrteLUT[4195] = 16'hbb37;
RsqrteLUT[4196] = 16'hbb33;
RsqrteLUT[4197] = 16'hbb2f;
RsqrteLUT[4198] = 16'hbb2b;
RsqrteLUT[4199] = 16'hbb27;
RsqrteLUT[4200] = 16'hbb23;
RsqrteLUT[4201] = 16'hbb1f;
RsqrteLUT[4202] = 16'hbb1b;
RsqrteLUT[4203] = 16'hbb17;
RsqrteLUT[4204] = 16'hbb14;
RsqrteLUT[4205] = 16'hbb10;
RsqrteLUT[4206] = 16'hbb0d;
RsqrteLUT[4207] = 16'hbb09;
RsqrteLUT[4208] = 16'hbb06;
RsqrteLUT[4209] = 16'hbb02;
RsqrteLUT[4210] = 16'hbaff;
RsqrteLUT[4211] = 16'hbafb;
RsqrteLUT[4212] = 16'hbaf8;
RsqrteLUT[4213] = 16'hbaf5;
RsqrteLUT[4214] = 16'hbaf2;
RsqrteLUT[4215] = 16'hbaee;
RsqrteLUT[4216] = 16'hbaeb;
RsqrteLUT[4217] = 16'hbae8;
RsqrteLUT[4218] = 16'hbae5;
RsqrteLUT[4219] = 16'hbae2;
RsqrteLUT[4220] = 16'hbadf;
RsqrteLUT[4221] = 16'hbadc;
RsqrteLUT[4222] = 16'hbad9;
RsqrteLUT[4223] = 16'hbad6;
RsqrteLUT[4224] = 16'hbad4;
RsqrteLUT[4225] = 16'hbace;
RsqrteLUT[4226] = 16'hbac9;
RsqrteLUT[4227] = 16'hbac3;
RsqrteLUT[4228] = 16'hbabe;
RsqrteLUT[4229] = 16'hbab9;
RsqrteLUT[4230] = 16'hbab4;
RsqrteLUT[4231] = 16'hbaaf;
RsqrteLUT[4232] = 16'hbaaa;
RsqrteLUT[4233] = 16'hbaa5;
RsqrteLUT[4234] = 16'hbaa1;
RsqrteLUT[4235] = 16'hba9c;
RsqrteLUT[4236] = 16'hba98;
RsqrteLUT[4237] = 16'hba94;
RsqrteLUT[4238] = 16'hba8f;
RsqrteLUT[4239] = 16'hba8b;
RsqrteLUT[4240] = 16'hba87;
RsqrteLUT[4241] = 16'hba83;
RsqrteLUT[4242] = 16'hba7f;
RsqrteLUT[4243] = 16'hba7b;
RsqrteLUT[4244] = 16'hba78;
RsqrteLUT[4245] = 16'hba74;
RsqrteLUT[4246] = 16'hba70;
RsqrteLUT[4247] = 16'hba6d;
RsqrteLUT[4248] = 16'hba69;
RsqrteLUT[4249] = 16'hba66;
RsqrteLUT[4250] = 16'hba62;
RsqrteLUT[4251] = 16'hba5f;
RsqrteLUT[4252] = 16'hba5b;
RsqrteLUT[4253] = 16'hba58;
RsqrteLUT[4254] = 16'hba55;
RsqrteLUT[4255] = 16'hba52;
RsqrteLUT[4256] = 16'hba4f;
RsqrteLUT[4257] = 16'hba4c;
RsqrteLUT[4258] = 16'hba49;
RsqrteLUT[4259] = 16'hba46;
RsqrteLUT[4260] = 16'hba43;
RsqrteLUT[4261] = 16'hba40;
RsqrteLUT[4262] = 16'hba3d;
RsqrteLUT[4263] = 16'hba3a;
RsqrteLUT[4264] = 16'hba38;
RsqrteLUT[4265] = 16'hba35;
RsqrteLUT[4266] = 16'hba32;
RsqrteLUT[4267] = 16'hba2f;
RsqrteLUT[4268] = 16'hba2d;
RsqrteLUT[4269] = 16'hba2a;
RsqrteLUT[4270] = 16'hba28;
RsqrteLUT[4271] = 16'hba25;
RsqrteLUT[4272] = 16'hba23;
RsqrteLUT[4273] = 16'hba20;
RsqrteLUT[4274] = 16'hba1e;
RsqrteLUT[4275] = 16'hba1c;
RsqrteLUT[4276] = 16'hba19;
RsqrteLUT[4277] = 16'hba17;
RsqrteLUT[4278] = 16'hba15;
RsqrteLUT[4279] = 16'hba13;
RsqrteLUT[4280] = 16'hba10;
RsqrteLUT[4281] = 16'hba0e;
RsqrteLUT[4282] = 16'hba0c;
RsqrteLUT[4283] = 16'hba0a;
RsqrteLUT[4284] = 16'hba08;
RsqrteLUT[4285] = 16'hba06;
RsqrteLUT[4286] = 16'hba04;
RsqrteLUT[4287] = 16'hba02;
RsqrteLUT[4288] = 16'hba00;
RsqrteLUT[4289] = 16'hb9f8;
RsqrteLUT[4290] = 16'hb9f0;
RsqrteLUT[4291] = 16'hb9e8;
RsqrteLUT[4292] = 16'hb9e1;
RsqrteLUT[4293] = 16'hb9da;
RsqrteLUT[4294] = 16'hb9d3;
RsqrteLUT[4295] = 16'hb9cc;
RsqrteLUT[4296] = 16'hb9c5;
RsqrteLUT[4297] = 16'hb9be;
RsqrteLUT[4298] = 16'hb9b8;
RsqrteLUT[4299] = 16'hb9b1;
RsqrteLUT[4300] = 16'hb9ab;
RsqrteLUT[4301] = 16'hb9a5;
RsqrteLUT[4302] = 16'hb99f;
RsqrteLUT[4303] = 16'hb999;
RsqrteLUT[4304] = 16'hb993;
RsqrteLUT[4305] = 16'hb98e;
RsqrteLUT[4306] = 16'hb988;
RsqrteLUT[4307] = 16'hb983;
RsqrteLUT[4308] = 16'hb97d;
RsqrteLUT[4309] = 16'hb978;
RsqrteLUT[4310] = 16'hb973;
RsqrteLUT[4311] = 16'hb96e;
RsqrteLUT[4312] = 16'hb969;
RsqrteLUT[4313] = 16'hb964;
RsqrteLUT[4314] = 16'hb95f;
RsqrteLUT[4315] = 16'hb95a;
RsqrteLUT[4316] = 16'hb956;
RsqrteLUT[4317] = 16'hb951;
RsqrteLUT[4318] = 16'hb94c;
RsqrteLUT[4319] = 16'hb948;
RsqrteLUT[4320] = 16'hb944;
RsqrteLUT[4321] = 16'hb93f;
RsqrteLUT[4322] = 16'hb93b;
RsqrteLUT[4323] = 16'hb937;
RsqrteLUT[4324] = 16'hb933;
RsqrteLUT[4325] = 16'hb92f;
RsqrteLUT[4326] = 16'hb92b;
RsqrteLUT[4327] = 16'hb927;
RsqrteLUT[4328] = 16'hb923;
RsqrteLUT[4329] = 16'hb91f;
RsqrteLUT[4330] = 16'hb91b;
RsqrteLUT[4331] = 16'hb917;
RsqrteLUT[4332] = 16'hb914;
RsqrteLUT[4333] = 16'hb910;
RsqrteLUT[4334] = 16'hb90d;
RsqrteLUT[4335] = 16'hb909;
RsqrteLUT[4336] = 16'hb906;
RsqrteLUT[4337] = 16'hb902;
RsqrteLUT[4338] = 16'hb8ff;
RsqrteLUT[4339] = 16'hb8fb;
RsqrteLUT[4340] = 16'hb8f8;
RsqrteLUT[4341] = 16'hb8f5;
RsqrteLUT[4342] = 16'hb8f2;
RsqrteLUT[4343] = 16'hb8ee;
RsqrteLUT[4344] = 16'hb8eb;
RsqrteLUT[4345] = 16'hb8e8;
RsqrteLUT[4346] = 16'hb8e5;
RsqrteLUT[4347] = 16'hb8e2;
RsqrteLUT[4348] = 16'hb8df;
RsqrteLUT[4349] = 16'hb8dc;
RsqrteLUT[4350] = 16'hb8d9;
RsqrteLUT[4351] = 16'hb8d6;
RsqrteLUT[4352] = 16'hb8d4;
RsqrteLUT[4353] = 16'hb8ce;
RsqrteLUT[4354] = 16'hb8c9;
RsqrteLUT[4355] = 16'hb8c3;
RsqrteLUT[4356] = 16'hb8be;
RsqrteLUT[4357] = 16'hb8b9;
RsqrteLUT[4358] = 16'hb8b4;
RsqrteLUT[4359] = 16'hb8af;
RsqrteLUT[4360] = 16'hb8aa;
RsqrteLUT[4361] = 16'hb8a5;
RsqrteLUT[4362] = 16'hb8a1;
RsqrteLUT[4363] = 16'hb89c;
RsqrteLUT[4364] = 16'hb898;
RsqrteLUT[4365] = 16'hb894;
RsqrteLUT[4366] = 16'hb88f;
RsqrteLUT[4367] = 16'hb88b;
RsqrteLUT[4368] = 16'hb887;
RsqrteLUT[4369] = 16'hb883;
RsqrteLUT[4370] = 16'hb87f;
RsqrteLUT[4371] = 16'hb87b;
RsqrteLUT[4372] = 16'hb878;
RsqrteLUT[4373] = 16'hb874;
RsqrteLUT[4374] = 16'hb870;
RsqrteLUT[4375] = 16'hb86d;
RsqrteLUT[4376] = 16'hb869;
RsqrteLUT[4377] = 16'hb866;
RsqrteLUT[4378] = 16'hb862;
RsqrteLUT[4379] = 16'hb85f;
RsqrteLUT[4380] = 16'hb85b;
RsqrteLUT[4381] = 16'hb858;
RsqrteLUT[4382] = 16'hb855;
RsqrteLUT[4383] = 16'hb852;
RsqrteLUT[4384] = 16'hb84f;
RsqrteLUT[4385] = 16'hb84c;
RsqrteLUT[4386] = 16'hb849;
RsqrteLUT[4387] = 16'hb846;
RsqrteLUT[4388] = 16'hb843;
RsqrteLUT[4389] = 16'hb840;
RsqrteLUT[4390] = 16'hb83d;
RsqrteLUT[4391] = 16'hb83a;
RsqrteLUT[4392] = 16'hb838;
RsqrteLUT[4393] = 16'hb835;
RsqrteLUT[4394] = 16'hb832;
RsqrteLUT[4395] = 16'hb82f;
RsqrteLUT[4396] = 16'hb82d;
RsqrteLUT[4397] = 16'hb82a;
RsqrteLUT[4398] = 16'hb828;
RsqrteLUT[4399] = 16'hb825;
RsqrteLUT[4400] = 16'hb823;
RsqrteLUT[4401] = 16'hb820;
RsqrteLUT[4402] = 16'hb81e;
RsqrteLUT[4403] = 16'hb81c;
RsqrteLUT[4404] = 16'hb819;
RsqrteLUT[4405] = 16'hb817;
RsqrteLUT[4406] = 16'hb815;
RsqrteLUT[4407] = 16'hb813;
RsqrteLUT[4408] = 16'hb810;
RsqrteLUT[4409] = 16'hb80e;
RsqrteLUT[4410] = 16'hb80c;
RsqrteLUT[4411] = 16'hb80a;
RsqrteLUT[4412] = 16'hb808;
RsqrteLUT[4413] = 16'hb806;
RsqrteLUT[4414] = 16'hb804;
RsqrteLUT[4415] = 16'hb802;
RsqrteLUT[4416] = 16'hb800;
RsqrteLUT[4417] = 16'hb7f8;
RsqrteLUT[4418] = 16'hb7f0;
RsqrteLUT[4419] = 16'hb7e8;
RsqrteLUT[4420] = 16'hb7e1;
RsqrteLUT[4421] = 16'hb7da;
RsqrteLUT[4422] = 16'hb7d3;
RsqrteLUT[4423] = 16'hb7cc;
RsqrteLUT[4424] = 16'hb7c5;
RsqrteLUT[4425] = 16'hb7be;
RsqrteLUT[4426] = 16'hb7b8;
RsqrteLUT[4427] = 16'hb7b1;
RsqrteLUT[4428] = 16'hb7ab;
RsqrteLUT[4429] = 16'hb7a5;
RsqrteLUT[4430] = 16'hb79f;
RsqrteLUT[4431] = 16'hb799;
RsqrteLUT[4432] = 16'hb793;
RsqrteLUT[4433] = 16'hb78e;
RsqrteLUT[4434] = 16'hb788;
RsqrteLUT[4435] = 16'hb783;
RsqrteLUT[4436] = 16'hb77d;
RsqrteLUT[4437] = 16'hb778;
RsqrteLUT[4438] = 16'hb773;
RsqrteLUT[4439] = 16'hb76e;
RsqrteLUT[4440] = 16'hb769;
RsqrteLUT[4441] = 16'hb764;
RsqrteLUT[4442] = 16'hb75f;
RsqrteLUT[4443] = 16'hb75a;
RsqrteLUT[4444] = 16'hb756;
RsqrteLUT[4445] = 16'hb751;
RsqrteLUT[4446] = 16'hb74c;
RsqrteLUT[4447] = 16'hb748;
RsqrteLUT[4448] = 16'hb744;
RsqrteLUT[4449] = 16'hb73f;
RsqrteLUT[4450] = 16'hb73b;
RsqrteLUT[4451] = 16'hb737;
RsqrteLUT[4452] = 16'hb733;
RsqrteLUT[4453] = 16'hb72f;
RsqrteLUT[4454] = 16'hb72b;
RsqrteLUT[4455] = 16'hb727;
RsqrteLUT[4456] = 16'hb723;
RsqrteLUT[4457] = 16'hb71f;
RsqrteLUT[4458] = 16'hb71b;
RsqrteLUT[4459] = 16'hb717;
RsqrteLUT[4460] = 16'hb714;
RsqrteLUT[4461] = 16'hb710;
RsqrteLUT[4462] = 16'hb70d;
RsqrteLUT[4463] = 16'hb709;
RsqrteLUT[4464] = 16'hb706;
RsqrteLUT[4465] = 16'hb702;
RsqrteLUT[4466] = 16'hb6ff;
RsqrteLUT[4467] = 16'hb6fb;
RsqrteLUT[4468] = 16'hb6f8;
RsqrteLUT[4469] = 16'hb6f5;
RsqrteLUT[4470] = 16'hb6f2;
RsqrteLUT[4471] = 16'hb6ee;
RsqrteLUT[4472] = 16'hb6eb;
RsqrteLUT[4473] = 16'hb6e8;
RsqrteLUT[4474] = 16'hb6e5;
RsqrteLUT[4475] = 16'hb6e2;
RsqrteLUT[4476] = 16'hb6df;
RsqrteLUT[4477] = 16'hb6dc;
RsqrteLUT[4478] = 16'hb6d9;
RsqrteLUT[4479] = 16'hb6d6;
RsqrteLUT[4480] = 16'hb6d4;
RsqrteLUT[4481] = 16'hb6ce;
RsqrteLUT[4482] = 16'hb6c9;
RsqrteLUT[4483] = 16'hb6c3;
RsqrteLUT[4484] = 16'hb6be;
RsqrteLUT[4485] = 16'hb6b9;
RsqrteLUT[4486] = 16'hb6b4;
RsqrteLUT[4487] = 16'hb6af;
RsqrteLUT[4488] = 16'hb6aa;
RsqrteLUT[4489] = 16'hb6a5;
RsqrteLUT[4490] = 16'hb6a1;
RsqrteLUT[4491] = 16'hb69c;
RsqrteLUT[4492] = 16'hb698;
RsqrteLUT[4493] = 16'hb694;
RsqrteLUT[4494] = 16'hb68f;
RsqrteLUT[4495] = 16'hb68b;
RsqrteLUT[4496] = 16'hb687;
RsqrteLUT[4497] = 16'hb683;
RsqrteLUT[4498] = 16'hb67f;
RsqrteLUT[4499] = 16'hb67b;
RsqrteLUT[4500] = 16'hb678;
RsqrteLUT[4501] = 16'hb674;
RsqrteLUT[4502] = 16'hb670;
RsqrteLUT[4503] = 16'hb66d;
RsqrteLUT[4504] = 16'hb669;
RsqrteLUT[4505] = 16'hb666;
RsqrteLUT[4506] = 16'hb662;
RsqrteLUT[4507] = 16'hb65f;
RsqrteLUT[4508] = 16'hb65b;
RsqrteLUT[4509] = 16'hb658;
RsqrteLUT[4510] = 16'hb655;
RsqrteLUT[4511] = 16'hb652;
RsqrteLUT[4512] = 16'hb64f;
RsqrteLUT[4513] = 16'hb64c;
RsqrteLUT[4514] = 16'hb649;
RsqrteLUT[4515] = 16'hb646;
RsqrteLUT[4516] = 16'hb643;
RsqrteLUT[4517] = 16'hb640;
RsqrteLUT[4518] = 16'hb63d;
RsqrteLUT[4519] = 16'hb63a;
RsqrteLUT[4520] = 16'hb638;
RsqrteLUT[4521] = 16'hb635;
RsqrteLUT[4522] = 16'hb632;
RsqrteLUT[4523] = 16'hb62f;
RsqrteLUT[4524] = 16'hb62d;
RsqrteLUT[4525] = 16'hb62a;
RsqrteLUT[4526] = 16'hb628;
RsqrteLUT[4527] = 16'hb625;
RsqrteLUT[4528] = 16'hb623;
RsqrteLUT[4529] = 16'hb620;
RsqrteLUT[4530] = 16'hb61e;
RsqrteLUT[4531] = 16'hb61c;
RsqrteLUT[4532] = 16'hb619;
RsqrteLUT[4533] = 16'hb617;
RsqrteLUT[4534] = 16'hb615;
RsqrteLUT[4535] = 16'hb613;
RsqrteLUT[4536] = 16'hb610;
RsqrteLUT[4537] = 16'hb60e;
RsqrteLUT[4538] = 16'hb60c;
RsqrteLUT[4539] = 16'hb60a;
RsqrteLUT[4540] = 16'hb608;
RsqrteLUT[4541] = 16'hb606;
RsqrteLUT[4542] = 16'hb604;
RsqrteLUT[4543] = 16'hb602;
RsqrteLUT[4544] = 16'hb600;
RsqrteLUT[4545] = 16'hb5f8;
RsqrteLUT[4546] = 16'hb5f0;
RsqrteLUT[4547] = 16'hb5e8;
RsqrteLUT[4548] = 16'hb5e1;
RsqrteLUT[4549] = 16'hb5da;
RsqrteLUT[4550] = 16'hb5d3;
RsqrteLUT[4551] = 16'hb5cc;
RsqrteLUT[4552] = 16'hb5c5;
RsqrteLUT[4553] = 16'hb5be;
RsqrteLUT[4554] = 16'hb5b8;
RsqrteLUT[4555] = 16'hb5b1;
RsqrteLUT[4556] = 16'hb5ab;
RsqrteLUT[4557] = 16'hb5a5;
RsqrteLUT[4558] = 16'hb59f;
RsqrteLUT[4559] = 16'hb599;
RsqrteLUT[4560] = 16'hb593;
RsqrteLUT[4561] = 16'hb58e;
RsqrteLUT[4562] = 16'hb588;
RsqrteLUT[4563] = 16'hb583;
RsqrteLUT[4564] = 16'hb57d;
RsqrteLUT[4565] = 16'hb578;
RsqrteLUT[4566] = 16'hb573;
RsqrteLUT[4567] = 16'hb56e;
RsqrteLUT[4568] = 16'hb569;
RsqrteLUT[4569] = 16'hb564;
RsqrteLUT[4570] = 16'hb55f;
RsqrteLUT[4571] = 16'hb55a;
RsqrteLUT[4572] = 16'hb556;
RsqrteLUT[4573] = 16'hb551;
RsqrteLUT[4574] = 16'hb54c;
RsqrteLUT[4575] = 16'hb548;
RsqrteLUT[4576] = 16'hb544;
RsqrteLUT[4577] = 16'hb53f;
RsqrteLUT[4578] = 16'hb53b;
RsqrteLUT[4579] = 16'hb537;
RsqrteLUT[4580] = 16'hb533;
RsqrteLUT[4581] = 16'hb52f;
RsqrteLUT[4582] = 16'hb52b;
RsqrteLUT[4583] = 16'hb527;
RsqrteLUT[4584] = 16'hb523;
RsqrteLUT[4585] = 16'hb51f;
RsqrteLUT[4586] = 16'hb51b;
RsqrteLUT[4587] = 16'hb517;
RsqrteLUT[4588] = 16'hb514;
RsqrteLUT[4589] = 16'hb510;
RsqrteLUT[4590] = 16'hb50d;
RsqrteLUT[4591] = 16'hb509;
RsqrteLUT[4592] = 16'hb506;
RsqrteLUT[4593] = 16'hb502;
RsqrteLUT[4594] = 16'hb4ff;
RsqrteLUT[4595] = 16'hb4fb;
RsqrteLUT[4596] = 16'hb4f8;
RsqrteLUT[4597] = 16'hb4f5;
RsqrteLUT[4598] = 16'hb4f2;
RsqrteLUT[4599] = 16'hb4ee;
RsqrteLUT[4600] = 16'hb4eb;
RsqrteLUT[4601] = 16'hb4e8;
RsqrteLUT[4602] = 16'hb4e5;
RsqrteLUT[4603] = 16'hb4e2;
RsqrteLUT[4604] = 16'hb4df;
RsqrteLUT[4605] = 16'hb4dc;
RsqrteLUT[4606] = 16'hb4d9;
RsqrteLUT[4607] = 16'hb4d6;
RsqrteLUT[4608] = 16'hb4d4;
RsqrteLUT[4609] = 16'hb4ce;
RsqrteLUT[4610] = 16'hb4c9;
RsqrteLUT[4611] = 16'hb4c3;
RsqrteLUT[4612] = 16'hb4be;
RsqrteLUT[4613] = 16'hb4b9;
RsqrteLUT[4614] = 16'hb4b4;
RsqrteLUT[4615] = 16'hb4af;
RsqrteLUT[4616] = 16'hb4aa;
RsqrteLUT[4617] = 16'hb4a5;
RsqrteLUT[4618] = 16'hb4a1;
RsqrteLUT[4619] = 16'hb49c;
RsqrteLUT[4620] = 16'hb498;
RsqrteLUT[4621] = 16'hb494;
RsqrteLUT[4622] = 16'hb48f;
RsqrteLUT[4623] = 16'hb48b;
RsqrteLUT[4624] = 16'hb487;
RsqrteLUT[4625] = 16'hb483;
RsqrteLUT[4626] = 16'hb47f;
RsqrteLUT[4627] = 16'hb47b;
RsqrteLUT[4628] = 16'hb478;
RsqrteLUT[4629] = 16'hb474;
RsqrteLUT[4630] = 16'hb470;
RsqrteLUT[4631] = 16'hb46d;
RsqrteLUT[4632] = 16'hb469;
RsqrteLUT[4633] = 16'hb466;
RsqrteLUT[4634] = 16'hb462;
RsqrteLUT[4635] = 16'hb45f;
RsqrteLUT[4636] = 16'hb45b;
RsqrteLUT[4637] = 16'hb458;
RsqrteLUT[4638] = 16'hb455;
RsqrteLUT[4639] = 16'hb452;
RsqrteLUT[4640] = 16'hb44f;
RsqrteLUT[4641] = 16'hb44c;
RsqrteLUT[4642] = 16'hb449;
RsqrteLUT[4643] = 16'hb446;
RsqrteLUT[4644] = 16'hb443;
RsqrteLUT[4645] = 16'hb440;
RsqrteLUT[4646] = 16'hb43d;
RsqrteLUT[4647] = 16'hb43a;
RsqrteLUT[4648] = 16'hb438;
RsqrteLUT[4649] = 16'hb435;
RsqrteLUT[4650] = 16'hb432;
RsqrteLUT[4651] = 16'hb42f;
RsqrteLUT[4652] = 16'hb42d;
RsqrteLUT[4653] = 16'hb42a;
RsqrteLUT[4654] = 16'hb428;
RsqrteLUT[4655] = 16'hb425;
RsqrteLUT[4656] = 16'hb423;
RsqrteLUT[4657] = 16'hb420;
RsqrteLUT[4658] = 16'hb41e;
RsqrteLUT[4659] = 16'hb41c;
RsqrteLUT[4660] = 16'hb419;
RsqrteLUT[4661] = 16'hb417;
RsqrteLUT[4662] = 16'hb415;
RsqrteLUT[4663] = 16'hb413;
RsqrteLUT[4664] = 16'hb410;
RsqrteLUT[4665] = 16'hb40e;
RsqrteLUT[4666] = 16'hb40c;
RsqrteLUT[4667] = 16'hb40a;
RsqrteLUT[4668] = 16'hb408;
RsqrteLUT[4669] = 16'hb406;
RsqrteLUT[4670] = 16'hb404;
RsqrteLUT[4671] = 16'hb402;
RsqrteLUT[4672] = 16'hb400;
RsqrteLUT[4673] = 16'hb3f8;
RsqrteLUT[4674] = 16'hb3f0;
RsqrteLUT[4675] = 16'hb3e8;
RsqrteLUT[4676] = 16'hb3e1;
RsqrteLUT[4677] = 16'hb3da;
RsqrteLUT[4678] = 16'hb3d3;
RsqrteLUT[4679] = 16'hb3cc;
RsqrteLUT[4680] = 16'hb3c5;
RsqrteLUT[4681] = 16'hb3be;
RsqrteLUT[4682] = 16'hb3b8;
RsqrteLUT[4683] = 16'hb3b1;
RsqrteLUT[4684] = 16'hb3ab;
RsqrteLUT[4685] = 16'hb3a5;
RsqrteLUT[4686] = 16'hb39f;
RsqrteLUT[4687] = 16'hb399;
RsqrteLUT[4688] = 16'hb393;
RsqrteLUT[4689] = 16'hb38e;
RsqrteLUT[4690] = 16'hb388;
RsqrteLUT[4691] = 16'hb383;
RsqrteLUT[4692] = 16'hb37d;
RsqrteLUT[4693] = 16'hb378;
RsqrteLUT[4694] = 16'hb373;
RsqrteLUT[4695] = 16'hb36e;
RsqrteLUT[4696] = 16'hb369;
RsqrteLUT[4697] = 16'hb364;
RsqrteLUT[4698] = 16'hb35f;
RsqrteLUT[4699] = 16'hb35a;
RsqrteLUT[4700] = 16'hb356;
RsqrteLUT[4701] = 16'hb351;
RsqrteLUT[4702] = 16'hb34c;
RsqrteLUT[4703] = 16'hb348;
RsqrteLUT[4704] = 16'hb344;
RsqrteLUT[4705] = 16'hb33f;
RsqrteLUT[4706] = 16'hb33b;
RsqrteLUT[4707] = 16'hb337;
RsqrteLUT[4708] = 16'hb333;
RsqrteLUT[4709] = 16'hb32f;
RsqrteLUT[4710] = 16'hb32b;
RsqrteLUT[4711] = 16'hb327;
RsqrteLUT[4712] = 16'hb323;
RsqrteLUT[4713] = 16'hb31f;
RsqrteLUT[4714] = 16'hb31b;
RsqrteLUT[4715] = 16'hb317;
RsqrteLUT[4716] = 16'hb314;
RsqrteLUT[4717] = 16'hb310;
RsqrteLUT[4718] = 16'hb30d;
RsqrteLUT[4719] = 16'hb309;
RsqrteLUT[4720] = 16'hb306;
RsqrteLUT[4721] = 16'hb302;
RsqrteLUT[4722] = 16'hb2ff;
RsqrteLUT[4723] = 16'hb2fb;
RsqrteLUT[4724] = 16'hb2f8;
RsqrteLUT[4725] = 16'hb2f5;
RsqrteLUT[4726] = 16'hb2f2;
RsqrteLUT[4727] = 16'hb2ee;
RsqrteLUT[4728] = 16'hb2eb;
RsqrteLUT[4729] = 16'hb2e8;
RsqrteLUT[4730] = 16'hb2e5;
RsqrteLUT[4731] = 16'hb2e2;
RsqrteLUT[4732] = 16'hb2df;
RsqrteLUT[4733] = 16'hb2dc;
RsqrteLUT[4734] = 16'hb2d9;
RsqrteLUT[4735] = 16'hb2d6;
RsqrteLUT[4736] = 16'hb2d4;
RsqrteLUT[4737] = 16'hb2ce;
RsqrteLUT[4738] = 16'hb2c9;
RsqrteLUT[4739] = 16'hb2c3;
RsqrteLUT[4740] = 16'hb2be;
RsqrteLUT[4741] = 16'hb2b9;
RsqrteLUT[4742] = 16'hb2b4;
RsqrteLUT[4743] = 16'hb2af;
RsqrteLUT[4744] = 16'hb2aa;
RsqrteLUT[4745] = 16'hb2a5;
RsqrteLUT[4746] = 16'hb2a1;
RsqrteLUT[4747] = 16'hb29c;
RsqrteLUT[4748] = 16'hb298;
RsqrteLUT[4749] = 16'hb294;
RsqrteLUT[4750] = 16'hb28f;
RsqrteLUT[4751] = 16'hb28b;
RsqrteLUT[4752] = 16'hb287;
RsqrteLUT[4753] = 16'hb283;
RsqrteLUT[4754] = 16'hb27f;
RsqrteLUT[4755] = 16'hb27b;
RsqrteLUT[4756] = 16'hb278;
RsqrteLUT[4757] = 16'hb274;
RsqrteLUT[4758] = 16'hb270;
RsqrteLUT[4759] = 16'hb26d;
RsqrteLUT[4760] = 16'hb269;
RsqrteLUT[4761] = 16'hb266;
RsqrteLUT[4762] = 16'hb262;
RsqrteLUT[4763] = 16'hb25f;
RsqrteLUT[4764] = 16'hb25b;
RsqrteLUT[4765] = 16'hb258;
RsqrteLUT[4766] = 16'hb255;
RsqrteLUT[4767] = 16'hb252;
RsqrteLUT[4768] = 16'hb24f;
RsqrteLUT[4769] = 16'hb24c;
RsqrteLUT[4770] = 16'hb249;
RsqrteLUT[4771] = 16'hb246;
RsqrteLUT[4772] = 16'hb243;
RsqrteLUT[4773] = 16'hb240;
RsqrteLUT[4774] = 16'hb23d;
RsqrteLUT[4775] = 16'hb23a;
RsqrteLUT[4776] = 16'hb238;
RsqrteLUT[4777] = 16'hb235;
RsqrteLUT[4778] = 16'hb232;
RsqrteLUT[4779] = 16'hb22f;
RsqrteLUT[4780] = 16'hb22d;
RsqrteLUT[4781] = 16'hb22a;
RsqrteLUT[4782] = 16'hb228;
RsqrteLUT[4783] = 16'hb225;
RsqrteLUT[4784] = 16'hb223;
RsqrteLUT[4785] = 16'hb220;
RsqrteLUT[4786] = 16'hb21e;
RsqrteLUT[4787] = 16'hb21c;
RsqrteLUT[4788] = 16'hb219;
RsqrteLUT[4789] = 16'hb217;
RsqrteLUT[4790] = 16'hb215;
RsqrteLUT[4791] = 16'hb213;
RsqrteLUT[4792] = 16'hb210;
RsqrteLUT[4793] = 16'hb20e;
RsqrteLUT[4794] = 16'hb20c;
RsqrteLUT[4795] = 16'hb20a;
RsqrteLUT[4796] = 16'hb208;
RsqrteLUT[4797] = 16'hb206;
RsqrteLUT[4798] = 16'hb204;
RsqrteLUT[4799] = 16'hb202;
RsqrteLUT[4800] = 16'hb200;
RsqrteLUT[4801] = 16'hb1f8;
RsqrteLUT[4802] = 16'hb1f0;
RsqrteLUT[4803] = 16'hb1e8;
RsqrteLUT[4804] = 16'hb1e1;
RsqrteLUT[4805] = 16'hb1da;
RsqrteLUT[4806] = 16'hb1d3;
RsqrteLUT[4807] = 16'hb1cc;
RsqrteLUT[4808] = 16'hb1c5;
RsqrteLUT[4809] = 16'hb1be;
RsqrteLUT[4810] = 16'hb1b8;
RsqrteLUT[4811] = 16'hb1b1;
RsqrteLUT[4812] = 16'hb1ab;
RsqrteLUT[4813] = 16'hb1a5;
RsqrteLUT[4814] = 16'hb19f;
RsqrteLUT[4815] = 16'hb199;
RsqrteLUT[4816] = 16'hb193;
RsqrteLUT[4817] = 16'hb18e;
RsqrteLUT[4818] = 16'hb188;
RsqrteLUT[4819] = 16'hb183;
RsqrteLUT[4820] = 16'hb17d;
RsqrteLUT[4821] = 16'hb178;
RsqrteLUT[4822] = 16'hb173;
RsqrteLUT[4823] = 16'hb16e;
RsqrteLUT[4824] = 16'hb169;
RsqrteLUT[4825] = 16'hb164;
RsqrteLUT[4826] = 16'hb15f;
RsqrteLUT[4827] = 16'hb15a;
RsqrteLUT[4828] = 16'hb156;
RsqrteLUT[4829] = 16'hb151;
RsqrteLUT[4830] = 16'hb14c;
RsqrteLUT[4831] = 16'hb148;
RsqrteLUT[4832] = 16'hb144;
RsqrteLUT[4833] = 16'hb13f;
RsqrteLUT[4834] = 16'hb13b;
RsqrteLUT[4835] = 16'hb137;
RsqrteLUT[4836] = 16'hb133;
RsqrteLUT[4837] = 16'hb12f;
RsqrteLUT[4838] = 16'hb12b;
RsqrteLUT[4839] = 16'hb127;
RsqrteLUT[4840] = 16'hb123;
RsqrteLUT[4841] = 16'hb11f;
RsqrteLUT[4842] = 16'hb11b;
RsqrteLUT[4843] = 16'hb117;
RsqrteLUT[4844] = 16'hb114;
RsqrteLUT[4845] = 16'hb110;
RsqrteLUT[4846] = 16'hb10d;
RsqrteLUT[4847] = 16'hb109;
RsqrteLUT[4848] = 16'hb106;
RsqrteLUT[4849] = 16'hb102;
RsqrteLUT[4850] = 16'hb0ff;
RsqrteLUT[4851] = 16'hb0fb;
RsqrteLUT[4852] = 16'hb0f8;
RsqrteLUT[4853] = 16'hb0f5;
RsqrteLUT[4854] = 16'hb0f2;
RsqrteLUT[4855] = 16'hb0ee;
RsqrteLUT[4856] = 16'hb0eb;
RsqrteLUT[4857] = 16'hb0e8;
RsqrteLUT[4858] = 16'hb0e5;
RsqrteLUT[4859] = 16'hb0e2;
RsqrteLUT[4860] = 16'hb0df;
RsqrteLUT[4861] = 16'hb0dc;
RsqrteLUT[4862] = 16'hb0d9;
RsqrteLUT[4863] = 16'hb0d6;
RsqrteLUT[4864] = 16'hb0d4;
RsqrteLUT[4865] = 16'hb0ce;
RsqrteLUT[4866] = 16'hb0c9;
RsqrteLUT[4867] = 16'hb0c3;
RsqrteLUT[4868] = 16'hb0be;
RsqrteLUT[4869] = 16'hb0b9;
RsqrteLUT[4870] = 16'hb0b4;
RsqrteLUT[4871] = 16'hb0af;
RsqrteLUT[4872] = 16'hb0aa;
RsqrteLUT[4873] = 16'hb0a5;
RsqrteLUT[4874] = 16'hb0a1;
RsqrteLUT[4875] = 16'hb09c;
RsqrteLUT[4876] = 16'hb098;
RsqrteLUT[4877] = 16'hb094;
RsqrteLUT[4878] = 16'hb08f;
RsqrteLUT[4879] = 16'hb08b;
RsqrteLUT[4880] = 16'hb087;
RsqrteLUT[4881] = 16'hb083;
RsqrteLUT[4882] = 16'hb07f;
RsqrteLUT[4883] = 16'hb07b;
RsqrteLUT[4884] = 16'hb078;
RsqrteLUT[4885] = 16'hb074;
RsqrteLUT[4886] = 16'hb070;
RsqrteLUT[4887] = 16'hb06d;
RsqrteLUT[4888] = 16'hb069;
RsqrteLUT[4889] = 16'hb066;
RsqrteLUT[4890] = 16'hb062;
RsqrteLUT[4891] = 16'hb05f;
RsqrteLUT[4892] = 16'hb05b;
RsqrteLUT[4893] = 16'hb058;
RsqrteLUT[4894] = 16'hb055;
RsqrteLUT[4895] = 16'hb052;
RsqrteLUT[4896] = 16'hb04f;
RsqrteLUT[4897] = 16'hb04c;
RsqrteLUT[4898] = 16'hb049;
RsqrteLUT[4899] = 16'hb046;
RsqrteLUT[4900] = 16'hb043;
RsqrteLUT[4901] = 16'hb040;
RsqrteLUT[4902] = 16'hb03d;
RsqrteLUT[4903] = 16'hb03a;
RsqrteLUT[4904] = 16'hb038;
RsqrteLUT[4905] = 16'hb035;
RsqrteLUT[4906] = 16'hb032;
RsqrteLUT[4907] = 16'hb02f;
RsqrteLUT[4908] = 16'hb02d;
RsqrteLUT[4909] = 16'hb02a;
RsqrteLUT[4910] = 16'hb028;
RsqrteLUT[4911] = 16'hb025;
RsqrteLUT[4912] = 16'hb023;
RsqrteLUT[4913] = 16'hb020;
RsqrteLUT[4914] = 16'hb01e;
RsqrteLUT[4915] = 16'hb01c;
RsqrteLUT[4916] = 16'hb019;
RsqrteLUT[4917] = 16'hb017;
RsqrteLUT[4918] = 16'hb015;
RsqrteLUT[4919] = 16'hb013;
RsqrteLUT[4920] = 16'hb010;
RsqrteLUT[4921] = 16'hb00e;
RsqrteLUT[4922] = 16'hb00c;
RsqrteLUT[4923] = 16'hb00a;
RsqrteLUT[4924] = 16'hb008;
RsqrteLUT[4925] = 16'hb006;
RsqrteLUT[4926] = 16'hb004;
RsqrteLUT[4927] = 16'hb002;
RsqrteLUT[4928] = 16'hb000;
RsqrteLUT[4929] = 16'haff8;
RsqrteLUT[4930] = 16'haff0;
RsqrteLUT[4931] = 16'hafe8;
RsqrteLUT[4932] = 16'hafe1;
RsqrteLUT[4933] = 16'hafda;
RsqrteLUT[4934] = 16'hafd3;
RsqrteLUT[4935] = 16'hafcc;
RsqrteLUT[4936] = 16'hafc5;
RsqrteLUT[4937] = 16'hafbe;
RsqrteLUT[4938] = 16'hafb8;
RsqrteLUT[4939] = 16'hafb1;
RsqrteLUT[4940] = 16'hafab;
RsqrteLUT[4941] = 16'hafa5;
RsqrteLUT[4942] = 16'haf9f;
RsqrteLUT[4943] = 16'haf99;
RsqrteLUT[4944] = 16'haf93;
RsqrteLUT[4945] = 16'haf8e;
RsqrteLUT[4946] = 16'haf88;
RsqrteLUT[4947] = 16'haf83;
RsqrteLUT[4948] = 16'haf7d;
RsqrteLUT[4949] = 16'haf78;
RsqrteLUT[4950] = 16'haf73;
RsqrteLUT[4951] = 16'haf6e;
RsqrteLUT[4952] = 16'haf69;
RsqrteLUT[4953] = 16'haf64;
RsqrteLUT[4954] = 16'haf5f;
RsqrteLUT[4955] = 16'haf5a;
RsqrteLUT[4956] = 16'haf56;
RsqrteLUT[4957] = 16'haf51;
RsqrteLUT[4958] = 16'haf4c;
RsqrteLUT[4959] = 16'haf48;
RsqrteLUT[4960] = 16'haf44;
RsqrteLUT[4961] = 16'haf3f;
RsqrteLUT[4962] = 16'haf3b;
RsqrteLUT[4963] = 16'haf37;
RsqrteLUT[4964] = 16'haf33;
RsqrteLUT[4965] = 16'haf2f;
RsqrteLUT[4966] = 16'haf2b;
RsqrteLUT[4967] = 16'haf27;
RsqrteLUT[4968] = 16'haf23;
RsqrteLUT[4969] = 16'haf1f;
RsqrteLUT[4970] = 16'haf1b;
RsqrteLUT[4971] = 16'haf17;
RsqrteLUT[4972] = 16'haf14;
RsqrteLUT[4973] = 16'haf10;
RsqrteLUT[4974] = 16'haf0d;
RsqrteLUT[4975] = 16'haf09;
RsqrteLUT[4976] = 16'haf06;
RsqrteLUT[4977] = 16'haf02;
RsqrteLUT[4978] = 16'haeff;
RsqrteLUT[4979] = 16'haefb;
RsqrteLUT[4980] = 16'haef8;
RsqrteLUT[4981] = 16'haef5;
RsqrteLUT[4982] = 16'haef2;
RsqrteLUT[4983] = 16'haeee;
RsqrteLUT[4984] = 16'haeeb;
RsqrteLUT[4985] = 16'haee8;
RsqrteLUT[4986] = 16'haee5;
RsqrteLUT[4987] = 16'haee2;
RsqrteLUT[4988] = 16'haedf;
RsqrteLUT[4989] = 16'haedc;
RsqrteLUT[4990] = 16'haed9;
RsqrteLUT[4991] = 16'haed6;
RsqrteLUT[4992] = 16'haed4;
RsqrteLUT[4993] = 16'haece;
RsqrteLUT[4994] = 16'haec9;
RsqrteLUT[4995] = 16'haec3;
RsqrteLUT[4996] = 16'haebe;
RsqrteLUT[4997] = 16'haeb9;
RsqrteLUT[4998] = 16'haeb4;
RsqrteLUT[4999] = 16'haeaf;
RsqrteLUT[5000] = 16'haeaa;
RsqrteLUT[5001] = 16'haea5;
RsqrteLUT[5002] = 16'haea1;
RsqrteLUT[5003] = 16'hae9c;
RsqrteLUT[5004] = 16'hae98;
RsqrteLUT[5005] = 16'hae94;
RsqrteLUT[5006] = 16'hae8f;
RsqrteLUT[5007] = 16'hae8b;
RsqrteLUT[5008] = 16'hae87;
RsqrteLUT[5009] = 16'hae83;
RsqrteLUT[5010] = 16'hae7f;
RsqrteLUT[5011] = 16'hae7b;
RsqrteLUT[5012] = 16'hae78;
RsqrteLUT[5013] = 16'hae74;
RsqrteLUT[5014] = 16'hae70;
RsqrteLUT[5015] = 16'hae6d;
RsqrteLUT[5016] = 16'hae69;
RsqrteLUT[5017] = 16'hae66;
RsqrteLUT[5018] = 16'hae62;
RsqrteLUT[5019] = 16'hae5f;
RsqrteLUT[5020] = 16'hae5b;
RsqrteLUT[5021] = 16'hae58;
RsqrteLUT[5022] = 16'hae55;
RsqrteLUT[5023] = 16'hae52;
RsqrteLUT[5024] = 16'hae4f;
RsqrteLUT[5025] = 16'hae4c;
RsqrteLUT[5026] = 16'hae49;
RsqrteLUT[5027] = 16'hae46;
RsqrteLUT[5028] = 16'hae43;
RsqrteLUT[5029] = 16'hae40;
RsqrteLUT[5030] = 16'hae3d;
RsqrteLUT[5031] = 16'hae3a;
RsqrteLUT[5032] = 16'hae38;
RsqrteLUT[5033] = 16'hae35;
RsqrteLUT[5034] = 16'hae32;
RsqrteLUT[5035] = 16'hae2f;
RsqrteLUT[5036] = 16'hae2d;
RsqrteLUT[5037] = 16'hae2a;
RsqrteLUT[5038] = 16'hae28;
RsqrteLUT[5039] = 16'hae25;
RsqrteLUT[5040] = 16'hae23;
RsqrteLUT[5041] = 16'hae20;
RsqrteLUT[5042] = 16'hae1e;
RsqrteLUT[5043] = 16'hae1c;
RsqrteLUT[5044] = 16'hae19;
RsqrteLUT[5045] = 16'hae17;
RsqrteLUT[5046] = 16'hae15;
RsqrteLUT[5047] = 16'hae13;
RsqrteLUT[5048] = 16'hae10;
RsqrteLUT[5049] = 16'hae0e;
RsqrteLUT[5050] = 16'hae0c;
RsqrteLUT[5051] = 16'hae0a;
RsqrteLUT[5052] = 16'hae08;
RsqrteLUT[5053] = 16'hae06;
RsqrteLUT[5054] = 16'hae04;
RsqrteLUT[5055] = 16'hae02;
RsqrteLUT[5056] = 16'hae00;
RsqrteLUT[5057] = 16'hadf8;
RsqrteLUT[5058] = 16'hadf0;
RsqrteLUT[5059] = 16'hade8;
RsqrteLUT[5060] = 16'hade1;
RsqrteLUT[5061] = 16'hadda;
RsqrteLUT[5062] = 16'hadd3;
RsqrteLUT[5063] = 16'hadcc;
RsqrteLUT[5064] = 16'hadc5;
RsqrteLUT[5065] = 16'hadbe;
RsqrteLUT[5066] = 16'hadb8;
RsqrteLUT[5067] = 16'hadb1;
RsqrteLUT[5068] = 16'hadab;
RsqrteLUT[5069] = 16'hada5;
RsqrteLUT[5070] = 16'had9f;
RsqrteLUT[5071] = 16'had99;
RsqrteLUT[5072] = 16'had93;
RsqrteLUT[5073] = 16'had8e;
RsqrteLUT[5074] = 16'had88;
RsqrteLUT[5075] = 16'had83;
RsqrteLUT[5076] = 16'had7d;
RsqrteLUT[5077] = 16'had78;
RsqrteLUT[5078] = 16'had73;
RsqrteLUT[5079] = 16'had6e;
RsqrteLUT[5080] = 16'had69;
RsqrteLUT[5081] = 16'had64;
RsqrteLUT[5082] = 16'had5f;
RsqrteLUT[5083] = 16'had5a;
RsqrteLUT[5084] = 16'had56;
RsqrteLUT[5085] = 16'had51;
RsqrteLUT[5086] = 16'had4c;
RsqrteLUT[5087] = 16'had48;
RsqrteLUT[5088] = 16'had44;
RsqrteLUT[5089] = 16'had3f;
RsqrteLUT[5090] = 16'had3b;
RsqrteLUT[5091] = 16'had37;
RsqrteLUT[5092] = 16'had33;
RsqrteLUT[5093] = 16'had2f;
RsqrteLUT[5094] = 16'had2b;
RsqrteLUT[5095] = 16'had27;
RsqrteLUT[5096] = 16'had23;
RsqrteLUT[5097] = 16'had1f;
RsqrteLUT[5098] = 16'had1b;
RsqrteLUT[5099] = 16'had17;
RsqrteLUT[5100] = 16'had14;
RsqrteLUT[5101] = 16'had10;
RsqrteLUT[5102] = 16'had0d;
RsqrteLUT[5103] = 16'had09;
RsqrteLUT[5104] = 16'had06;
RsqrteLUT[5105] = 16'had02;
RsqrteLUT[5106] = 16'hacff;
RsqrteLUT[5107] = 16'hacfb;
RsqrteLUT[5108] = 16'hacf8;
RsqrteLUT[5109] = 16'hacf5;
RsqrteLUT[5110] = 16'hacf2;
RsqrteLUT[5111] = 16'hacee;
RsqrteLUT[5112] = 16'haceb;
RsqrteLUT[5113] = 16'hace8;
RsqrteLUT[5114] = 16'hace5;
RsqrteLUT[5115] = 16'hace2;
RsqrteLUT[5116] = 16'hacdf;
RsqrteLUT[5117] = 16'hacdc;
RsqrteLUT[5118] = 16'hacd9;
RsqrteLUT[5119] = 16'hacd6;
RsqrteLUT[5120] = 16'hacd4;
RsqrteLUT[5121] = 16'hacce;
RsqrteLUT[5122] = 16'hacc9;
RsqrteLUT[5123] = 16'hacc3;
RsqrteLUT[5124] = 16'hacbe;
RsqrteLUT[5125] = 16'hacb9;
RsqrteLUT[5126] = 16'hacb4;
RsqrteLUT[5127] = 16'hacaf;
RsqrteLUT[5128] = 16'hacaa;
RsqrteLUT[5129] = 16'haca5;
RsqrteLUT[5130] = 16'haca1;
RsqrteLUT[5131] = 16'hac9c;
RsqrteLUT[5132] = 16'hac98;
RsqrteLUT[5133] = 16'hac94;
RsqrteLUT[5134] = 16'hac8f;
RsqrteLUT[5135] = 16'hac8b;
RsqrteLUT[5136] = 16'hac87;
RsqrteLUT[5137] = 16'hac83;
RsqrteLUT[5138] = 16'hac7f;
RsqrteLUT[5139] = 16'hac7b;
RsqrteLUT[5140] = 16'hac78;
RsqrteLUT[5141] = 16'hac74;
RsqrteLUT[5142] = 16'hac70;
RsqrteLUT[5143] = 16'hac6d;
RsqrteLUT[5144] = 16'hac69;
RsqrteLUT[5145] = 16'hac66;
RsqrteLUT[5146] = 16'hac62;
RsqrteLUT[5147] = 16'hac5f;
RsqrteLUT[5148] = 16'hac5b;
RsqrteLUT[5149] = 16'hac58;
RsqrteLUT[5150] = 16'hac55;
RsqrteLUT[5151] = 16'hac52;
RsqrteLUT[5152] = 16'hac4f;
RsqrteLUT[5153] = 16'hac4c;
RsqrteLUT[5154] = 16'hac49;
RsqrteLUT[5155] = 16'hac46;
RsqrteLUT[5156] = 16'hac43;
RsqrteLUT[5157] = 16'hac40;
RsqrteLUT[5158] = 16'hac3d;
RsqrteLUT[5159] = 16'hac3a;
RsqrteLUT[5160] = 16'hac38;
RsqrteLUT[5161] = 16'hac35;
RsqrteLUT[5162] = 16'hac32;
RsqrteLUT[5163] = 16'hac2f;
RsqrteLUT[5164] = 16'hac2d;
RsqrteLUT[5165] = 16'hac2a;
RsqrteLUT[5166] = 16'hac28;
RsqrteLUT[5167] = 16'hac25;
RsqrteLUT[5168] = 16'hac23;
RsqrteLUT[5169] = 16'hac20;
RsqrteLUT[5170] = 16'hac1e;
RsqrteLUT[5171] = 16'hac1c;
RsqrteLUT[5172] = 16'hac19;
RsqrteLUT[5173] = 16'hac17;
RsqrteLUT[5174] = 16'hac15;
RsqrteLUT[5175] = 16'hac13;
RsqrteLUT[5176] = 16'hac10;
RsqrteLUT[5177] = 16'hac0e;
RsqrteLUT[5178] = 16'hac0c;
RsqrteLUT[5179] = 16'hac0a;
RsqrteLUT[5180] = 16'hac08;
RsqrteLUT[5181] = 16'hac06;
RsqrteLUT[5182] = 16'hac04;
RsqrteLUT[5183] = 16'hac02;
RsqrteLUT[5184] = 16'hac00;
RsqrteLUT[5185] = 16'habf8;
RsqrteLUT[5186] = 16'habf0;
RsqrteLUT[5187] = 16'habe8;
RsqrteLUT[5188] = 16'habe1;
RsqrteLUT[5189] = 16'habda;
RsqrteLUT[5190] = 16'habd3;
RsqrteLUT[5191] = 16'habcc;
RsqrteLUT[5192] = 16'habc5;
RsqrteLUT[5193] = 16'habbe;
RsqrteLUT[5194] = 16'habb8;
RsqrteLUT[5195] = 16'habb1;
RsqrteLUT[5196] = 16'habab;
RsqrteLUT[5197] = 16'haba5;
RsqrteLUT[5198] = 16'hab9f;
RsqrteLUT[5199] = 16'hab99;
RsqrteLUT[5200] = 16'hab93;
RsqrteLUT[5201] = 16'hab8e;
RsqrteLUT[5202] = 16'hab88;
RsqrteLUT[5203] = 16'hab83;
RsqrteLUT[5204] = 16'hab7d;
RsqrteLUT[5205] = 16'hab78;
RsqrteLUT[5206] = 16'hab73;
RsqrteLUT[5207] = 16'hab6e;
RsqrteLUT[5208] = 16'hab69;
RsqrteLUT[5209] = 16'hab64;
RsqrteLUT[5210] = 16'hab5f;
RsqrteLUT[5211] = 16'hab5a;
RsqrteLUT[5212] = 16'hab56;
RsqrteLUT[5213] = 16'hab51;
RsqrteLUT[5214] = 16'hab4c;
RsqrteLUT[5215] = 16'hab48;
RsqrteLUT[5216] = 16'hab44;
RsqrteLUT[5217] = 16'hab3f;
RsqrteLUT[5218] = 16'hab3b;
RsqrteLUT[5219] = 16'hab37;
RsqrteLUT[5220] = 16'hab33;
RsqrteLUT[5221] = 16'hab2f;
RsqrteLUT[5222] = 16'hab2b;
RsqrteLUT[5223] = 16'hab27;
RsqrteLUT[5224] = 16'hab23;
RsqrteLUT[5225] = 16'hab1f;
RsqrteLUT[5226] = 16'hab1b;
RsqrteLUT[5227] = 16'hab17;
RsqrteLUT[5228] = 16'hab14;
RsqrteLUT[5229] = 16'hab10;
RsqrteLUT[5230] = 16'hab0d;
RsqrteLUT[5231] = 16'hab09;
RsqrteLUT[5232] = 16'hab06;
RsqrteLUT[5233] = 16'hab02;
RsqrteLUT[5234] = 16'haaff;
RsqrteLUT[5235] = 16'haafb;
RsqrteLUT[5236] = 16'haaf8;
RsqrteLUT[5237] = 16'haaf5;
RsqrteLUT[5238] = 16'haaf2;
RsqrteLUT[5239] = 16'haaee;
RsqrteLUT[5240] = 16'haaeb;
RsqrteLUT[5241] = 16'haae8;
RsqrteLUT[5242] = 16'haae5;
RsqrteLUT[5243] = 16'haae2;
RsqrteLUT[5244] = 16'haadf;
RsqrteLUT[5245] = 16'haadc;
RsqrteLUT[5246] = 16'haad9;
RsqrteLUT[5247] = 16'haad6;
RsqrteLUT[5248] = 16'haad4;
RsqrteLUT[5249] = 16'haace;
RsqrteLUT[5250] = 16'haac9;
RsqrteLUT[5251] = 16'haac3;
RsqrteLUT[5252] = 16'haabe;
RsqrteLUT[5253] = 16'haab9;
RsqrteLUT[5254] = 16'haab4;
RsqrteLUT[5255] = 16'haaaf;
RsqrteLUT[5256] = 16'haaaa;
RsqrteLUT[5257] = 16'haaa5;
RsqrteLUT[5258] = 16'haaa1;
RsqrteLUT[5259] = 16'haa9c;
RsqrteLUT[5260] = 16'haa98;
RsqrteLUT[5261] = 16'haa94;
RsqrteLUT[5262] = 16'haa8f;
RsqrteLUT[5263] = 16'haa8b;
RsqrteLUT[5264] = 16'haa87;
RsqrteLUT[5265] = 16'haa83;
RsqrteLUT[5266] = 16'haa7f;
RsqrteLUT[5267] = 16'haa7b;
RsqrteLUT[5268] = 16'haa78;
RsqrteLUT[5269] = 16'haa74;
RsqrteLUT[5270] = 16'haa70;
RsqrteLUT[5271] = 16'haa6d;
RsqrteLUT[5272] = 16'haa69;
RsqrteLUT[5273] = 16'haa66;
RsqrteLUT[5274] = 16'haa62;
RsqrteLUT[5275] = 16'haa5f;
RsqrteLUT[5276] = 16'haa5b;
RsqrteLUT[5277] = 16'haa58;
RsqrteLUT[5278] = 16'haa55;
RsqrteLUT[5279] = 16'haa52;
RsqrteLUT[5280] = 16'haa4f;
RsqrteLUT[5281] = 16'haa4c;
RsqrteLUT[5282] = 16'haa49;
RsqrteLUT[5283] = 16'haa46;
RsqrteLUT[5284] = 16'haa43;
RsqrteLUT[5285] = 16'haa40;
RsqrteLUT[5286] = 16'haa3d;
RsqrteLUT[5287] = 16'haa3a;
RsqrteLUT[5288] = 16'haa38;
RsqrteLUT[5289] = 16'haa35;
RsqrteLUT[5290] = 16'haa32;
RsqrteLUT[5291] = 16'haa2f;
RsqrteLUT[5292] = 16'haa2d;
RsqrteLUT[5293] = 16'haa2a;
RsqrteLUT[5294] = 16'haa28;
RsqrteLUT[5295] = 16'haa25;
RsqrteLUT[5296] = 16'haa23;
RsqrteLUT[5297] = 16'haa20;
RsqrteLUT[5298] = 16'haa1e;
RsqrteLUT[5299] = 16'haa1c;
RsqrteLUT[5300] = 16'haa19;
RsqrteLUT[5301] = 16'haa17;
RsqrteLUT[5302] = 16'haa15;
RsqrteLUT[5303] = 16'haa13;
RsqrteLUT[5304] = 16'haa10;
RsqrteLUT[5305] = 16'haa0e;
RsqrteLUT[5306] = 16'haa0c;
RsqrteLUT[5307] = 16'haa0a;
RsqrteLUT[5308] = 16'haa08;
RsqrteLUT[5309] = 16'haa06;
RsqrteLUT[5310] = 16'haa04;
RsqrteLUT[5311] = 16'haa02;
RsqrteLUT[5312] = 16'haa00;
RsqrteLUT[5313] = 16'ha9f8;
RsqrteLUT[5314] = 16'ha9f0;
RsqrteLUT[5315] = 16'ha9e8;
RsqrteLUT[5316] = 16'ha9e1;
RsqrteLUT[5317] = 16'ha9da;
RsqrteLUT[5318] = 16'ha9d3;
RsqrteLUT[5319] = 16'ha9cc;
RsqrteLUT[5320] = 16'ha9c5;
RsqrteLUT[5321] = 16'ha9be;
RsqrteLUT[5322] = 16'ha9b8;
RsqrteLUT[5323] = 16'ha9b1;
RsqrteLUT[5324] = 16'ha9ab;
RsqrteLUT[5325] = 16'ha9a5;
RsqrteLUT[5326] = 16'ha99f;
RsqrteLUT[5327] = 16'ha999;
RsqrteLUT[5328] = 16'ha993;
RsqrteLUT[5329] = 16'ha98e;
RsqrteLUT[5330] = 16'ha988;
RsqrteLUT[5331] = 16'ha983;
RsqrteLUT[5332] = 16'ha97d;
RsqrteLUT[5333] = 16'ha978;
RsqrteLUT[5334] = 16'ha973;
RsqrteLUT[5335] = 16'ha96e;
RsqrteLUT[5336] = 16'ha969;
RsqrteLUT[5337] = 16'ha964;
RsqrteLUT[5338] = 16'ha95f;
RsqrteLUT[5339] = 16'ha95a;
RsqrteLUT[5340] = 16'ha956;
RsqrteLUT[5341] = 16'ha951;
RsqrteLUT[5342] = 16'ha94c;
RsqrteLUT[5343] = 16'ha948;
RsqrteLUT[5344] = 16'ha944;
RsqrteLUT[5345] = 16'ha93f;
RsqrteLUT[5346] = 16'ha93b;
RsqrteLUT[5347] = 16'ha937;
RsqrteLUT[5348] = 16'ha933;
RsqrteLUT[5349] = 16'ha92f;
RsqrteLUT[5350] = 16'ha92b;
RsqrteLUT[5351] = 16'ha927;
RsqrteLUT[5352] = 16'ha923;
RsqrteLUT[5353] = 16'ha91f;
RsqrteLUT[5354] = 16'ha91b;
RsqrteLUT[5355] = 16'ha917;
RsqrteLUT[5356] = 16'ha914;
RsqrteLUT[5357] = 16'ha910;
RsqrteLUT[5358] = 16'ha90d;
RsqrteLUT[5359] = 16'ha909;
RsqrteLUT[5360] = 16'ha906;
RsqrteLUT[5361] = 16'ha902;
RsqrteLUT[5362] = 16'ha8ff;
RsqrteLUT[5363] = 16'ha8fb;
RsqrteLUT[5364] = 16'ha8f8;
RsqrteLUT[5365] = 16'ha8f5;
RsqrteLUT[5366] = 16'ha8f2;
RsqrteLUT[5367] = 16'ha8ee;
RsqrteLUT[5368] = 16'ha8eb;
RsqrteLUT[5369] = 16'ha8e8;
RsqrteLUT[5370] = 16'ha8e5;
RsqrteLUT[5371] = 16'ha8e2;
RsqrteLUT[5372] = 16'ha8df;
RsqrteLUT[5373] = 16'ha8dc;
RsqrteLUT[5374] = 16'ha8d9;
RsqrteLUT[5375] = 16'ha8d6;
RsqrteLUT[5376] = 16'ha8d4;
RsqrteLUT[5377] = 16'ha8ce;
RsqrteLUT[5378] = 16'ha8c9;
RsqrteLUT[5379] = 16'ha8c3;
RsqrteLUT[5380] = 16'ha8be;
RsqrteLUT[5381] = 16'ha8b9;
RsqrteLUT[5382] = 16'ha8b4;
RsqrteLUT[5383] = 16'ha8af;
RsqrteLUT[5384] = 16'ha8aa;
RsqrteLUT[5385] = 16'ha8a5;
RsqrteLUT[5386] = 16'ha8a1;
RsqrteLUT[5387] = 16'ha89c;
RsqrteLUT[5388] = 16'ha898;
RsqrteLUT[5389] = 16'ha894;
RsqrteLUT[5390] = 16'ha88f;
RsqrteLUT[5391] = 16'ha88b;
RsqrteLUT[5392] = 16'ha887;
RsqrteLUT[5393] = 16'ha883;
RsqrteLUT[5394] = 16'ha87f;
RsqrteLUT[5395] = 16'ha87b;
RsqrteLUT[5396] = 16'ha878;
RsqrteLUT[5397] = 16'ha874;
RsqrteLUT[5398] = 16'ha870;
RsqrteLUT[5399] = 16'ha86d;
RsqrteLUT[5400] = 16'ha869;
RsqrteLUT[5401] = 16'ha866;
RsqrteLUT[5402] = 16'ha862;
RsqrteLUT[5403] = 16'ha85f;
RsqrteLUT[5404] = 16'ha85b;
RsqrteLUT[5405] = 16'ha858;
RsqrteLUT[5406] = 16'ha855;
RsqrteLUT[5407] = 16'ha852;
RsqrteLUT[5408] = 16'ha84f;
RsqrteLUT[5409] = 16'ha84c;
RsqrteLUT[5410] = 16'ha849;
RsqrteLUT[5411] = 16'ha846;
RsqrteLUT[5412] = 16'ha843;
RsqrteLUT[5413] = 16'ha840;
RsqrteLUT[5414] = 16'ha83d;
RsqrteLUT[5415] = 16'ha83a;
RsqrteLUT[5416] = 16'ha838;
RsqrteLUT[5417] = 16'ha835;
RsqrteLUT[5418] = 16'ha832;
RsqrteLUT[5419] = 16'ha82f;
RsqrteLUT[5420] = 16'ha82d;
RsqrteLUT[5421] = 16'ha82a;
RsqrteLUT[5422] = 16'ha828;
RsqrteLUT[5423] = 16'ha825;
RsqrteLUT[5424] = 16'ha823;
RsqrteLUT[5425] = 16'ha820;
RsqrteLUT[5426] = 16'ha81e;
RsqrteLUT[5427] = 16'ha81c;
RsqrteLUT[5428] = 16'ha819;
RsqrteLUT[5429] = 16'ha817;
RsqrteLUT[5430] = 16'ha815;
RsqrteLUT[5431] = 16'ha813;
RsqrteLUT[5432] = 16'ha810;
RsqrteLUT[5433] = 16'ha80e;
RsqrteLUT[5434] = 16'ha80c;
RsqrteLUT[5435] = 16'ha80a;
RsqrteLUT[5436] = 16'ha808;
RsqrteLUT[5437] = 16'ha806;
RsqrteLUT[5438] = 16'ha804;
RsqrteLUT[5439] = 16'ha802;
RsqrteLUT[5440] = 16'ha800;
RsqrteLUT[5441] = 16'ha7f8;
RsqrteLUT[5442] = 16'ha7f0;
RsqrteLUT[5443] = 16'ha7e8;
RsqrteLUT[5444] = 16'ha7e1;
RsqrteLUT[5445] = 16'ha7da;
RsqrteLUT[5446] = 16'ha7d3;
RsqrteLUT[5447] = 16'ha7cc;
RsqrteLUT[5448] = 16'ha7c5;
RsqrteLUT[5449] = 16'ha7be;
RsqrteLUT[5450] = 16'ha7b8;
RsqrteLUT[5451] = 16'ha7b1;
RsqrteLUT[5452] = 16'ha7ab;
RsqrteLUT[5453] = 16'ha7a5;
RsqrteLUT[5454] = 16'ha79f;
RsqrteLUT[5455] = 16'ha799;
RsqrteLUT[5456] = 16'ha793;
RsqrteLUT[5457] = 16'ha78e;
RsqrteLUT[5458] = 16'ha788;
RsqrteLUT[5459] = 16'ha783;
RsqrteLUT[5460] = 16'ha77d;
RsqrteLUT[5461] = 16'ha778;
RsqrteLUT[5462] = 16'ha773;
RsqrteLUT[5463] = 16'ha76e;
RsqrteLUT[5464] = 16'ha769;
RsqrteLUT[5465] = 16'ha764;
RsqrteLUT[5466] = 16'ha75f;
RsqrteLUT[5467] = 16'ha75a;
RsqrteLUT[5468] = 16'ha756;
RsqrteLUT[5469] = 16'ha751;
RsqrteLUT[5470] = 16'ha74c;
RsqrteLUT[5471] = 16'ha748;
RsqrteLUT[5472] = 16'ha744;
RsqrteLUT[5473] = 16'ha73f;
RsqrteLUT[5474] = 16'ha73b;
RsqrteLUT[5475] = 16'ha737;
RsqrteLUT[5476] = 16'ha733;
RsqrteLUT[5477] = 16'ha72f;
RsqrteLUT[5478] = 16'ha72b;
RsqrteLUT[5479] = 16'ha727;
RsqrteLUT[5480] = 16'ha723;
RsqrteLUT[5481] = 16'ha71f;
RsqrteLUT[5482] = 16'ha71b;
RsqrteLUT[5483] = 16'ha717;
RsqrteLUT[5484] = 16'ha714;
RsqrteLUT[5485] = 16'ha710;
RsqrteLUT[5486] = 16'ha70d;
RsqrteLUT[5487] = 16'ha709;
RsqrteLUT[5488] = 16'ha706;
RsqrteLUT[5489] = 16'ha702;
RsqrteLUT[5490] = 16'ha6ff;
RsqrteLUT[5491] = 16'ha6fb;
RsqrteLUT[5492] = 16'ha6f8;
RsqrteLUT[5493] = 16'ha6f5;
RsqrteLUT[5494] = 16'ha6f2;
RsqrteLUT[5495] = 16'ha6ee;
RsqrteLUT[5496] = 16'ha6eb;
RsqrteLUT[5497] = 16'ha6e8;
RsqrteLUT[5498] = 16'ha6e5;
RsqrteLUT[5499] = 16'ha6e2;
RsqrteLUT[5500] = 16'ha6df;
RsqrteLUT[5501] = 16'ha6dc;
RsqrteLUT[5502] = 16'ha6d9;
RsqrteLUT[5503] = 16'ha6d6;
RsqrteLUT[5504] = 16'ha6d4;
RsqrteLUT[5505] = 16'ha6ce;
RsqrteLUT[5506] = 16'ha6c9;
RsqrteLUT[5507] = 16'ha6c3;
RsqrteLUT[5508] = 16'ha6be;
RsqrteLUT[5509] = 16'ha6b9;
RsqrteLUT[5510] = 16'ha6b4;
RsqrteLUT[5511] = 16'ha6af;
RsqrteLUT[5512] = 16'ha6aa;
RsqrteLUT[5513] = 16'ha6a5;
RsqrteLUT[5514] = 16'ha6a1;
RsqrteLUT[5515] = 16'ha69c;
RsqrteLUT[5516] = 16'ha698;
RsqrteLUT[5517] = 16'ha694;
RsqrteLUT[5518] = 16'ha68f;
RsqrteLUT[5519] = 16'ha68b;
RsqrteLUT[5520] = 16'ha687;
RsqrteLUT[5521] = 16'ha683;
RsqrteLUT[5522] = 16'ha67f;
RsqrteLUT[5523] = 16'ha67b;
RsqrteLUT[5524] = 16'ha678;
RsqrteLUT[5525] = 16'ha674;
RsqrteLUT[5526] = 16'ha670;
RsqrteLUT[5527] = 16'ha66d;
RsqrteLUT[5528] = 16'ha669;
RsqrteLUT[5529] = 16'ha666;
RsqrteLUT[5530] = 16'ha662;
RsqrteLUT[5531] = 16'ha65f;
RsqrteLUT[5532] = 16'ha65b;
RsqrteLUT[5533] = 16'ha658;
RsqrteLUT[5534] = 16'ha655;
RsqrteLUT[5535] = 16'ha652;
RsqrteLUT[5536] = 16'ha64f;
RsqrteLUT[5537] = 16'ha64c;
RsqrteLUT[5538] = 16'ha649;
RsqrteLUT[5539] = 16'ha646;
RsqrteLUT[5540] = 16'ha643;
RsqrteLUT[5541] = 16'ha640;
RsqrteLUT[5542] = 16'ha63d;
RsqrteLUT[5543] = 16'ha63a;
RsqrteLUT[5544] = 16'ha638;
RsqrteLUT[5545] = 16'ha635;
RsqrteLUT[5546] = 16'ha632;
RsqrteLUT[5547] = 16'ha62f;
RsqrteLUT[5548] = 16'ha62d;
RsqrteLUT[5549] = 16'ha62a;
RsqrteLUT[5550] = 16'ha628;
RsqrteLUT[5551] = 16'ha625;
RsqrteLUT[5552] = 16'ha623;
RsqrteLUT[5553] = 16'ha620;
RsqrteLUT[5554] = 16'ha61e;
RsqrteLUT[5555] = 16'ha61c;
RsqrteLUT[5556] = 16'ha619;
RsqrteLUT[5557] = 16'ha617;
RsqrteLUT[5558] = 16'ha615;
RsqrteLUT[5559] = 16'ha613;
RsqrteLUT[5560] = 16'ha610;
RsqrteLUT[5561] = 16'ha60e;
RsqrteLUT[5562] = 16'ha60c;
RsqrteLUT[5563] = 16'ha60a;
RsqrteLUT[5564] = 16'ha608;
RsqrteLUT[5565] = 16'ha606;
RsqrteLUT[5566] = 16'ha604;
RsqrteLUT[5567] = 16'ha602;
RsqrteLUT[5568] = 16'ha600;
RsqrteLUT[5569] = 16'ha5f8;
RsqrteLUT[5570] = 16'ha5f0;
RsqrteLUT[5571] = 16'ha5e8;
RsqrteLUT[5572] = 16'ha5e1;
RsqrteLUT[5573] = 16'ha5da;
RsqrteLUT[5574] = 16'ha5d3;
RsqrteLUT[5575] = 16'ha5cc;
RsqrteLUT[5576] = 16'ha5c5;
RsqrteLUT[5577] = 16'ha5be;
RsqrteLUT[5578] = 16'ha5b8;
RsqrteLUT[5579] = 16'ha5b1;
RsqrteLUT[5580] = 16'ha5ab;
RsqrteLUT[5581] = 16'ha5a5;
RsqrteLUT[5582] = 16'ha59f;
RsqrteLUT[5583] = 16'ha599;
RsqrteLUT[5584] = 16'ha593;
RsqrteLUT[5585] = 16'ha58e;
RsqrteLUT[5586] = 16'ha588;
RsqrteLUT[5587] = 16'ha583;
RsqrteLUT[5588] = 16'ha57d;
RsqrteLUT[5589] = 16'ha578;
RsqrteLUT[5590] = 16'ha573;
RsqrteLUT[5591] = 16'ha56e;
RsqrteLUT[5592] = 16'ha569;
RsqrteLUT[5593] = 16'ha564;
RsqrteLUT[5594] = 16'ha55f;
RsqrteLUT[5595] = 16'ha55a;
RsqrteLUT[5596] = 16'ha556;
RsqrteLUT[5597] = 16'ha551;
RsqrteLUT[5598] = 16'ha54c;
RsqrteLUT[5599] = 16'ha548;
RsqrteLUT[5600] = 16'ha544;
RsqrteLUT[5601] = 16'ha53f;
RsqrteLUT[5602] = 16'ha53b;
RsqrteLUT[5603] = 16'ha537;
RsqrteLUT[5604] = 16'ha533;
RsqrteLUT[5605] = 16'ha52f;
RsqrteLUT[5606] = 16'ha52b;
RsqrteLUT[5607] = 16'ha527;
RsqrteLUT[5608] = 16'ha523;
RsqrteLUT[5609] = 16'ha51f;
RsqrteLUT[5610] = 16'ha51b;
RsqrteLUT[5611] = 16'ha517;
RsqrteLUT[5612] = 16'ha514;
RsqrteLUT[5613] = 16'ha510;
RsqrteLUT[5614] = 16'ha50d;
RsqrteLUT[5615] = 16'ha509;
RsqrteLUT[5616] = 16'ha506;
RsqrteLUT[5617] = 16'ha502;
RsqrteLUT[5618] = 16'ha4ff;
RsqrteLUT[5619] = 16'ha4fb;
RsqrteLUT[5620] = 16'ha4f8;
RsqrteLUT[5621] = 16'ha4f5;
RsqrteLUT[5622] = 16'ha4f2;
RsqrteLUT[5623] = 16'ha4ee;
RsqrteLUT[5624] = 16'ha4eb;
RsqrteLUT[5625] = 16'ha4e8;
RsqrteLUT[5626] = 16'ha4e5;
RsqrteLUT[5627] = 16'ha4e2;
RsqrteLUT[5628] = 16'ha4df;
RsqrteLUT[5629] = 16'ha4dc;
RsqrteLUT[5630] = 16'ha4d9;
RsqrteLUT[5631] = 16'ha4d6;
RsqrteLUT[5632] = 16'ha4d4;
RsqrteLUT[5633] = 16'ha4ce;
RsqrteLUT[5634] = 16'ha4c9;
RsqrteLUT[5635] = 16'ha4c3;
RsqrteLUT[5636] = 16'ha4be;
RsqrteLUT[5637] = 16'ha4b9;
RsqrteLUT[5638] = 16'ha4b4;
RsqrteLUT[5639] = 16'ha4af;
RsqrteLUT[5640] = 16'ha4aa;
RsqrteLUT[5641] = 16'ha4a5;
RsqrteLUT[5642] = 16'ha4a1;
RsqrteLUT[5643] = 16'ha49c;
RsqrteLUT[5644] = 16'ha498;
RsqrteLUT[5645] = 16'ha494;
RsqrteLUT[5646] = 16'ha48f;
RsqrteLUT[5647] = 16'ha48b;
RsqrteLUT[5648] = 16'ha487;
RsqrteLUT[5649] = 16'ha483;
RsqrteLUT[5650] = 16'ha47f;
RsqrteLUT[5651] = 16'ha47b;
RsqrteLUT[5652] = 16'ha478;
RsqrteLUT[5653] = 16'ha474;
RsqrteLUT[5654] = 16'ha470;
RsqrteLUT[5655] = 16'ha46d;
RsqrteLUT[5656] = 16'ha469;
RsqrteLUT[5657] = 16'ha466;
RsqrteLUT[5658] = 16'ha462;
RsqrteLUT[5659] = 16'ha45f;
RsqrteLUT[5660] = 16'ha45b;
RsqrteLUT[5661] = 16'ha458;
RsqrteLUT[5662] = 16'ha455;
RsqrteLUT[5663] = 16'ha452;
RsqrteLUT[5664] = 16'ha44f;
RsqrteLUT[5665] = 16'ha44c;
RsqrteLUT[5666] = 16'ha449;
RsqrteLUT[5667] = 16'ha446;
RsqrteLUT[5668] = 16'ha443;
RsqrteLUT[5669] = 16'ha440;
RsqrteLUT[5670] = 16'ha43d;
RsqrteLUT[5671] = 16'ha43a;
RsqrteLUT[5672] = 16'ha438;
RsqrteLUT[5673] = 16'ha435;
RsqrteLUT[5674] = 16'ha432;
RsqrteLUT[5675] = 16'ha42f;
RsqrteLUT[5676] = 16'ha42d;
RsqrteLUT[5677] = 16'ha42a;
RsqrteLUT[5678] = 16'ha428;
RsqrteLUT[5679] = 16'ha425;
RsqrteLUT[5680] = 16'ha423;
RsqrteLUT[5681] = 16'ha420;
RsqrteLUT[5682] = 16'ha41e;
RsqrteLUT[5683] = 16'ha41c;
RsqrteLUT[5684] = 16'ha419;
RsqrteLUT[5685] = 16'ha417;
RsqrteLUT[5686] = 16'ha415;
RsqrteLUT[5687] = 16'ha413;
RsqrteLUT[5688] = 16'ha410;
RsqrteLUT[5689] = 16'ha40e;
RsqrteLUT[5690] = 16'ha40c;
RsqrteLUT[5691] = 16'ha40a;
RsqrteLUT[5692] = 16'ha408;
RsqrteLUT[5693] = 16'ha406;
RsqrteLUT[5694] = 16'ha404;
RsqrteLUT[5695] = 16'ha402;
RsqrteLUT[5696] = 16'ha400;
RsqrteLUT[5697] = 16'ha3f8;
RsqrteLUT[5698] = 16'ha3f0;
RsqrteLUT[5699] = 16'ha3e8;
RsqrteLUT[5700] = 16'ha3e1;
RsqrteLUT[5701] = 16'ha3da;
RsqrteLUT[5702] = 16'ha3d3;
RsqrteLUT[5703] = 16'ha3cc;
RsqrteLUT[5704] = 16'ha3c5;
RsqrteLUT[5705] = 16'ha3be;
RsqrteLUT[5706] = 16'ha3b8;
RsqrteLUT[5707] = 16'ha3b1;
RsqrteLUT[5708] = 16'ha3ab;
RsqrteLUT[5709] = 16'ha3a5;
RsqrteLUT[5710] = 16'ha39f;
RsqrteLUT[5711] = 16'ha399;
RsqrteLUT[5712] = 16'ha393;
RsqrteLUT[5713] = 16'ha38e;
RsqrteLUT[5714] = 16'ha388;
RsqrteLUT[5715] = 16'ha383;
RsqrteLUT[5716] = 16'ha37d;
RsqrteLUT[5717] = 16'ha378;
RsqrteLUT[5718] = 16'ha373;
RsqrteLUT[5719] = 16'ha36e;
RsqrteLUT[5720] = 16'ha369;
RsqrteLUT[5721] = 16'ha364;
RsqrteLUT[5722] = 16'ha35f;
RsqrteLUT[5723] = 16'ha35a;
RsqrteLUT[5724] = 16'ha356;
RsqrteLUT[5725] = 16'ha351;
RsqrteLUT[5726] = 16'ha34c;
RsqrteLUT[5727] = 16'ha348;
RsqrteLUT[5728] = 16'ha344;
RsqrteLUT[5729] = 16'ha33f;
RsqrteLUT[5730] = 16'ha33b;
RsqrteLUT[5731] = 16'ha337;
RsqrteLUT[5732] = 16'ha333;
RsqrteLUT[5733] = 16'ha32f;
RsqrteLUT[5734] = 16'ha32b;
RsqrteLUT[5735] = 16'ha327;
RsqrteLUT[5736] = 16'ha323;
RsqrteLUT[5737] = 16'ha31f;
RsqrteLUT[5738] = 16'ha31b;
RsqrteLUT[5739] = 16'ha317;
RsqrteLUT[5740] = 16'ha314;
RsqrteLUT[5741] = 16'ha310;
RsqrteLUT[5742] = 16'ha30d;
RsqrteLUT[5743] = 16'ha309;
RsqrteLUT[5744] = 16'ha306;
RsqrteLUT[5745] = 16'ha302;
RsqrteLUT[5746] = 16'ha2ff;
RsqrteLUT[5747] = 16'ha2fb;
RsqrteLUT[5748] = 16'ha2f8;
RsqrteLUT[5749] = 16'ha2f5;
RsqrteLUT[5750] = 16'ha2f2;
RsqrteLUT[5751] = 16'ha2ee;
RsqrteLUT[5752] = 16'ha2eb;
RsqrteLUT[5753] = 16'ha2e8;
RsqrteLUT[5754] = 16'ha2e5;
RsqrteLUT[5755] = 16'ha2e2;
RsqrteLUT[5756] = 16'ha2df;
RsqrteLUT[5757] = 16'ha2dc;
RsqrteLUT[5758] = 16'ha2d9;
RsqrteLUT[5759] = 16'ha2d6;
RsqrteLUT[5760] = 16'ha2d4;
RsqrteLUT[5761] = 16'ha2ce;
RsqrteLUT[5762] = 16'ha2c9;
RsqrteLUT[5763] = 16'ha2c3;
RsqrteLUT[5764] = 16'ha2be;
RsqrteLUT[5765] = 16'ha2b9;
RsqrteLUT[5766] = 16'ha2b4;
RsqrteLUT[5767] = 16'ha2af;
RsqrteLUT[5768] = 16'ha2aa;
RsqrteLUT[5769] = 16'ha2a5;
RsqrteLUT[5770] = 16'ha2a1;
RsqrteLUT[5771] = 16'ha29c;
RsqrteLUT[5772] = 16'ha298;
RsqrteLUT[5773] = 16'ha294;
RsqrteLUT[5774] = 16'ha28f;
RsqrteLUT[5775] = 16'ha28b;
RsqrteLUT[5776] = 16'ha287;
RsqrteLUT[5777] = 16'ha283;
RsqrteLUT[5778] = 16'ha27f;
RsqrteLUT[5779] = 16'ha27b;
RsqrteLUT[5780] = 16'ha278;
RsqrteLUT[5781] = 16'ha274;
RsqrteLUT[5782] = 16'ha270;
RsqrteLUT[5783] = 16'ha26d;
RsqrteLUT[5784] = 16'ha269;
RsqrteLUT[5785] = 16'ha266;
RsqrteLUT[5786] = 16'ha262;
RsqrteLUT[5787] = 16'ha25f;
RsqrteLUT[5788] = 16'ha25b;
RsqrteLUT[5789] = 16'ha258;
RsqrteLUT[5790] = 16'ha255;
RsqrteLUT[5791] = 16'ha252;
RsqrteLUT[5792] = 16'ha24f;
RsqrteLUT[5793] = 16'ha24c;
RsqrteLUT[5794] = 16'ha249;
RsqrteLUT[5795] = 16'ha246;
RsqrteLUT[5796] = 16'ha243;
RsqrteLUT[5797] = 16'ha240;
RsqrteLUT[5798] = 16'ha23d;
RsqrteLUT[5799] = 16'ha23a;
RsqrteLUT[5800] = 16'ha238;
RsqrteLUT[5801] = 16'ha235;
RsqrteLUT[5802] = 16'ha232;
RsqrteLUT[5803] = 16'ha22f;
RsqrteLUT[5804] = 16'ha22d;
RsqrteLUT[5805] = 16'ha22a;
RsqrteLUT[5806] = 16'ha228;
RsqrteLUT[5807] = 16'ha225;
RsqrteLUT[5808] = 16'ha223;
RsqrteLUT[5809] = 16'ha220;
RsqrteLUT[5810] = 16'ha21e;
RsqrteLUT[5811] = 16'ha21c;
RsqrteLUT[5812] = 16'ha219;
RsqrteLUT[5813] = 16'ha217;
RsqrteLUT[5814] = 16'ha215;
RsqrteLUT[5815] = 16'ha213;
RsqrteLUT[5816] = 16'ha210;
RsqrteLUT[5817] = 16'ha20e;
RsqrteLUT[5818] = 16'ha20c;
RsqrteLUT[5819] = 16'ha20a;
RsqrteLUT[5820] = 16'ha208;
RsqrteLUT[5821] = 16'ha206;
RsqrteLUT[5822] = 16'ha204;
RsqrteLUT[5823] = 16'ha202;
RsqrteLUT[5824] = 16'ha200;
RsqrteLUT[5825] = 16'ha1f8;
RsqrteLUT[5826] = 16'ha1f0;
RsqrteLUT[5827] = 16'ha1e8;
RsqrteLUT[5828] = 16'ha1e1;
RsqrteLUT[5829] = 16'ha1da;
RsqrteLUT[5830] = 16'ha1d3;
RsqrteLUT[5831] = 16'ha1cc;
RsqrteLUT[5832] = 16'ha1c5;
RsqrteLUT[5833] = 16'ha1be;
RsqrteLUT[5834] = 16'ha1b8;
RsqrteLUT[5835] = 16'ha1b1;
RsqrteLUT[5836] = 16'ha1ab;
RsqrteLUT[5837] = 16'ha1a5;
RsqrteLUT[5838] = 16'ha19f;
RsqrteLUT[5839] = 16'ha199;
RsqrteLUT[5840] = 16'ha193;
RsqrteLUT[5841] = 16'ha18e;
RsqrteLUT[5842] = 16'ha188;
RsqrteLUT[5843] = 16'ha183;
RsqrteLUT[5844] = 16'ha17d;
RsqrteLUT[5845] = 16'ha178;
RsqrteLUT[5846] = 16'ha173;
RsqrteLUT[5847] = 16'ha16e;
RsqrteLUT[5848] = 16'ha169;
RsqrteLUT[5849] = 16'ha164;
RsqrteLUT[5850] = 16'ha15f;
RsqrteLUT[5851] = 16'ha15a;
RsqrteLUT[5852] = 16'ha156;
RsqrteLUT[5853] = 16'ha151;
RsqrteLUT[5854] = 16'ha14c;
RsqrteLUT[5855] = 16'ha148;
RsqrteLUT[5856] = 16'ha144;
RsqrteLUT[5857] = 16'ha13f;
RsqrteLUT[5858] = 16'ha13b;
RsqrteLUT[5859] = 16'ha137;
RsqrteLUT[5860] = 16'ha133;
RsqrteLUT[5861] = 16'ha12f;
RsqrteLUT[5862] = 16'ha12b;
RsqrteLUT[5863] = 16'ha127;
RsqrteLUT[5864] = 16'ha123;
RsqrteLUT[5865] = 16'ha11f;
RsqrteLUT[5866] = 16'ha11b;
RsqrteLUT[5867] = 16'ha117;
RsqrteLUT[5868] = 16'ha114;
RsqrteLUT[5869] = 16'ha110;
RsqrteLUT[5870] = 16'ha10d;
RsqrteLUT[5871] = 16'ha109;
RsqrteLUT[5872] = 16'ha106;
RsqrteLUT[5873] = 16'ha102;
RsqrteLUT[5874] = 16'ha0ff;
RsqrteLUT[5875] = 16'ha0fb;
RsqrteLUT[5876] = 16'ha0f8;
RsqrteLUT[5877] = 16'ha0f5;
RsqrteLUT[5878] = 16'ha0f2;
RsqrteLUT[5879] = 16'ha0ee;
RsqrteLUT[5880] = 16'ha0eb;
RsqrteLUT[5881] = 16'ha0e8;
RsqrteLUT[5882] = 16'ha0e5;
RsqrteLUT[5883] = 16'ha0e2;
RsqrteLUT[5884] = 16'ha0df;
RsqrteLUT[5885] = 16'ha0dc;
RsqrteLUT[5886] = 16'ha0d9;
RsqrteLUT[5887] = 16'ha0d6;
RsqrteLUT[5888] = 16'ha0d4;
RsqrteLUT[5889] = 16'ha0ce;
RsqrteLUT[5890] = 16'ha0c9;
RsqrteLUT[5891] = 16'ha0c3;
RsqrteLUT[5892] = 16'ha0be;
RsqrteLUT[5893] = 16'ha0b9;
RsqrteLUT[5894] = 16'ha0b4;
RsqrteLUT[5895] = 16'ha0af;
RsqrteLUT[5896] = 16'ha0aa;
RsqrteLUT[5897] = 16'ha0a5;
RsqrteLUT[5898] = 16'ha0a1;
RsqrteLUT[5899] = 16'ha09c;
RsqrteLUT[5900] = 16'ha098;
RsqrteLUT[5901] = 16'ha094;
RsqrteLUT[5902] = 16'ha08f;
RsqrteLUT[5903] = 16'ha08b;
RsqrteLUT[5904] = 16'ha087;
RsqrteLUT[5905] = 16'ha083;
RsqrteLUT[5906] = 16'ha07f;
RsqrteLUT[5907] = 16'ha07b;
RsqrteLUT[5908] = 16'ha078;
RsqrteLUT[5909] = 16'ha074;
RsqrteLUT[5910] = 16'ha070;
RsqrteLUT[5911] = 16'ha06d;
RsqrteLUT[5912] = 16'ha069;
RsqrteLUT[5913] = 16'ha066;
RsqrteLUT[5914] = 16'ha062;
RsqrteLUT[5915] = 16'ha05f;
RsqrteLUT[5916] = 16'ha05b;
RsqrteLUT[5917] = 16'ha058;
RsqrteLUT[5918] = 16'ha055;
RsqrteLUT[5919] = 16'ha052;
RsqrteLUT[5920] = 16'ha04f;
RsqrteLUT[5921] = 16'ha04c;
RsqrteLUT[5922] = 16'ha049;
RsqrteLUT[5923] = 16'ha046;
RsqrteLUT[5924] = 16'ha043;
RsqrteLUT[5925] = 16'ha040;
RsqrteLUT[5926] = 16'ha03d;
RsqrteLUT[5927] = 16'ha03a;
RsqrteLUT[5928] = 16'ha038;
RsqrteLUT[5929] = 16'ha035;
RsqrteLUT[5930] = 16'ha032;
RsqrteLUT[5931] = 16'ha02f;
RsqrteLUT[5932] = 16'ha02d;
RsqrteLUT[5933] = 16'ha02a;
RsqrteLUT[5934] = 16'ha028;
RsqrteLUT[5935] = 16'ha025;
RsqrteLUT[5936] = 16'ha023;
RsqrteLUT[5937] = 16'ha020;
RsqrteLUT[5938] = 16'ha01e;
RsqrteLUT[5939] = 16'ha01c;
RsqrteLUT[5940] = 16'ha019;
RsqrteLUT[5941] = 16'ha017;
RsqrteLUT[5942] = 16'ha015;
RsqrteLUT[5943] = 16'ha013;
RsqrteLUT[5944] = 16'ha010;
RsqrteLUT[5945] = 16'ha00e;
RsqrteLUT[5946] = 16'ha00c;
RsqrteLUT[5947] = 16'ha00a;
RsqrteLUT[5948] = 16'ha008;
RsqrteLUT[5949] = 16'ha006;
RsqrteLUT[5950] = 16'ha004;
RsqrteLUT[5951] = 16'ha002;
RsqrteLUT[5952] = 16'ha000;
RsqrteLUT[5953] = 16'h9ff8;
RsqrteLUT[5954] = 16'h9ff0;
RsqrteLUT[5955] = 16'h9fe8;
RsqrteLUT[5956] = 16'h9fe1;
RsqrteLUT[5957] = 16'h9fda;
RsqrteLUT[5958] = 16'h9fd3;
RsqrteLUT[5959] = 16'h9fcc;
RsqrteLUT[5960] = 16'h9fc5;
RsqrteLUT[5961] = 16'h9fbe;
RsqrteLUT[5962] = 16'h9fb8;
RsqrteLUT[5963] = 16'h9fb1;
RsqrteLUT[5964] = 16'h9fab;
RsqrteLUT[5965] = 16'h9fa5;
RsqrteLUT[5966] = 16'h9f9f;
RsqrteLUT[5967] = 16'h9f99;
RsqrteLUT[5968] = 16'h9f93;
RsqrteLUT[5969] = 16'h9f8e;
RsqrteLUT[5970] = 16'h9f88;
RsqrteLUT[5971] = 16'h9f83;
RsqrteLUT[5972] = 16'h9f7d;
RsqrteLUT[5973] = 16'h9f78;
RsqrteLUT[5974] = 16'h9f73;
RsqrteLUT[5975] = 16'h9f6e;
RsqrteLUT[5976] = 16'h9f69;
RsqrteLUT[5977] = 16'h9f64;
RsqrteLUT[5978] = 16'h9f5f;
RsqrteLUT[5979] = 16'h9f5a;
RsqrteLUT[5980] = 16'h9f56;
RsqrteLUT[5981] = 16'h9f51;
RsqrteLUT[5982] = 16'h9f4c;
RsqrteLUT[5983] = 16'h9f48;
RsqrteLUT[5984] = 16'h9f44;
RsqrteLUT[5985] = 16'h9f3f;
RsqrteLUT[5986] = 16'h9f3b;
RsqrteLUT[5987] = 16'h9f37;
RsqrteLUT[5988] = 16'h9f33;
RsqrteLUT[5989] = 16'h9f2f;
RsqrteLUT[5990] = 16'h9f2b;
RsqrteLUT[5991] = 16'h9f27;
RsqrteLUT[5992] = 16'h9f23;
RsqrteLUT[5993] = 16'h9f1f;
RsqrteLUT[5994] = 16'h9f1b;
RsqrteLUT[5995] = 16'h9f17;
RsqrteLUT[5996] = 16'h9f14;
RsqrteLUT[5997] = 16'h9f10;
RsqrteLUT[5998] = 16'h9f0d;
RsqrteLUT[5999] = 16'h9f09;
RsqrteLUT[6000] = 16'h9f06;
RsqrteLUT[6001] = 16'h9f02;
RsqrteLUT[6002] = 16'h9eff;
RsqrteLUT[6003] = 16'h9efb;
RsqrteLUT[6004] = 16'h9ef8;
RsqrteLUT[6005] = 16'h9ef5;
RsqrteLUT[6006] = 16'h9ef2;
RsqrteLUT[6007] = 16'h9eee;
RsqrteLUT[6008] = 16'h9eeb;
RsqrteLUT[6009] = 16'h9ee8;
RsqrteLUT[6010] = 16'h9ee5;
RsqrteLUT[6011] = 16'h9ee2;
RsqrteLUT[6012] = 16'h9edf;
RsqrteLUT[6013] = 16'h9edc;
RsqrteLUT[6014] = 16'h9ed9;
RsqrteLUT[6015] = 16'h9ed6;
RsqrteLUT[6016] = 16'h9ed4;
RsqrteLUT[6017] = 16'h9ece;
RsqrteLUT[6018] = 16'h9ec9;
RsqrteLUT[6019] = 16'h9ec3;
RsqrteLUT[6020] = 16'h9ebe;
RsqrteLUT[6021] = 16'h9eb9;
RsqrteLUT[6022] = 16'h9eb4;
RsqrteLUT[6023] = 16'h9eaf;
RsqrteLUT[6024] = 16'h9eaa;
RsqrteLUT[6025] = 16'h9ea5;
RsqrteLUT[6026] = 16'h9ea1;
RsqrteLUT[6027] = 16'h9e9c;
RsqrteLUT[6028] = 16'h9e98;
RsqrteLUT[6029] = 16'h9e94;
RsqrteLUT[6030] = 16'h9e8f;
RsqrteLUT[6031] = 16'h9e8b;
RsqrteLUT[6032] = 16'h9e87;
RsqrteLUT[6033] = 16'h9e83;
RsqrteLUT[6034] = 16'h9e7f;
RsqrteLUT[6035] = 16'h9e7b;
RsqrteLUT[6036] = 16'h9e78;
RsqrteLUT[6037] = 16'h9e74;
RsqrteLUT[6038] = 16'h9e70;
RsqrteLUT[6039] = 16'h9e6d;
RsqrteLUT[6040] = 16'h9e69;
RsqrteLUT[6041] = 16'h9e66;
RsqrteLUT[6042] = 16'h9e62;
RsqrteLUT[6043] = 16'h9e5f;
RsqrteLUT[6044] = 16'h9e5b;
RsqrteLUT[6045] = 16'h9e58;
RsqrteLUT[6046] = 16'h9e55;
RsqrteLUT[6047] = 16'h9e52;
RsqrteLUT[6048] = 16'h9e4f;
RsqrteLUT[6049] = 16'h9e4c;
RsqrteLUT[6050] = 16'h9e49;
RsqrteLUT[6051] = 16'h9e46;
RsqrteLUT[6052] = 16'h9e43;
RsqrteLUT[6053] = 16'h9e40;
RsqrteLUT[6054] = 16'h9e3d;
RsqrteLUT[6055] = 16'h9e3a;
RsqrteLUT[6056] = 16'h9e38;
RsqrteLUT[6057] = 16'h9e35;
RsqrteLUT[6058] = 16'h9e32;
RsqrteLUT[6059] = 16'h9e2f;
RsqrteLUT[6060] = 16'h9e2d;
RsqrteLUT[6061] = 16'h9e2a;
RsqrteLUT[6062] = 16'h9e28;
RsqrteLUT[6063] = 16'h9e25;
RsqrteLUT[6064] = 16'h9e23;
RsqrteLUT[6065] = 16'h9e20;
RsqrteLUT[6066] = 16'h9e1e;
RsqrteLUT[6067] = 16'h9e1c;
RsqrteLUT[6068] = 16'h9e19;
RsqrteLUT[6069] = 16'h9e17;
RsqrteLUT[6070] = 16'h9e15;
RsqrteLUT[6071] = 16'h9e13;
RsqrteLUT[6072] = 16'h9e10;
RsqrteLUT[6073] = 16'h9e0e;
RsqrteLUT[6074] = 16'h9e0c;
RsqrteLUT[6075] = 16'h9e0a;
RsqrteLUT[6076] = 16'h9e08;
RsqrteLUT[6077] = 16'h9e06;
RsqrteLUT[6078] = 16'h9e04;
RsqrteLUT[6079] = 16'h9e02;
RsqrteLUT[6080] = 16'h9e00;
RsqrteLUT[6081] = 16'h9df8;
RsqrteLUT[6082] = 16'h9df0;
RsqrteLUT[6083] = 16'h9de8;
RsqrteLUT[6084] = 16'h9de1;
RsqrteLUT[6085] = 16'h9dda;
RsqrteLUT[6086] = 16'h9dd3;
RsqrteLUT[6087] = 16'h9dcc;
RsqrteLUT[6088] = 16'h9dc5;
RsqrteLUT[6089] = 16'h9dbe;
RsqrteLUT[6090] = 16'h9db8;
RsqrteLUT[6091] = 16'h9db1;
RsqrteLUT[6092] = 16'h9dab;
RsqrteLUT[6093] = 16'h9da5;
RsqrteLUT[6094] = 16'h9d9f;
RsqrteLUT[6095] = 16'h9d99;
RsqrteLUT[6096] = 16'h9d93;
RsqrteLUT[6097] = 16'h9d8e;
RsqrteLUT[6098] = 16'h9d88;
RsqrteLUT[6099] = 16'h9d83;
RsqrteLUT[6100] = 16'h9d7d;
RsqrteLUT[6101] = 16'h9d78;
RsqrteLUT[6102] = 16'h9d73;
RsqrteLUT[6103] = 16'h9d6e;
RsqrteLUT[6104] = 16'h9d69;
RsqrteLUT[6105] = 16'h9d64;
RsqrteLUT[6106] = 16'h9d5f;
RsqrteLUT[6107] = 16'h9d5a;
RsqrteLUT[6108] = 16'h9d56;
RsqrteLUT[6109] = 16'h9d51;
RsqrteLUT[6110] = 16'h9d4c;
RsqrteLUT[6111] = 16'h9d48;
RsqrteLUT[6112] = 16'h9d44;
RsqrteLUT[6113] = 16'h9d3f;
RsqrteLUT[6114] = 16'h9d3b;
RsqrteLUT[6115] = 16'h9d37;
RsqrteLUT[6116] = 16'h9d33;
RsqrteLUT[6117] = 16'h9d2f;
RsqrteLUT[6118] = 16'h9d2b;
RsqrteLUT[6119] = 16'h9d27;
RsqrteLUT[6120] = 16'h9d23;
RsqrteLUT[6121] = 16'h9d1f;
RsqrteLUT[6122] = 16'h9d1b;
RsqrteLUT[6123] = 16'h9d17;
RsqrteLUT[6124] = 16'h9d14;
RsqrteLUT[6125] = 16'h9d10;
RsqrteLUT[6126] = 16'h9d0d;
RsqrteLUT[6127] = 16'h9d09;
RsqrteLUT[6128] = 16'h9d06;
RsqrteLUT[6129] = 16'h9d02;
RsqrteLUT[6130] = 16'h9cff;
RsqrteLUT[6131] = 16'h9cfb;
RsqrteLUT[6132] = 16'h9cf8;
RsqrteLUT[6133] = 16'h9cf5;
RsqrteLUT[6134] = 16'h9cf2;
RsqrteLUT[6135] = 16'h9cee;
RsqrteLUT[6136] = 16'h9ceb;
RsqrteLUT[6137] = 16'h9ce8;
RsqrteLUT[6138] = 16'h9ce5;
RsqrteLUT[6139] = 16'h9ce2;
RsqrteLUT[6140] = 16'h9cdf;
RsqrteLUT[6141] = 16'h9cdc;
RsqrteLUT[6142] = 16'h9cd9;
RsqrteLUT[6143] = 16'h9cd6;
RsqrteLUT[6144] = 16'h9cd4;
RsqrteLUT[6145] = 16'h9cce;
RsqrteLUT[6146] = 16'h9cc9;
RsqrteLUT[6147] = 16'h9cc3;
RsqrteLUT[6148] = 16'h9cbe;
RsqrteLUT[6149] = 16'h9cb9;
RsqrteLUT[6150] = 16'h9cb4;
RsqrteLUT[6151] = 16'h9caf;
RsqrteLUT[6152] = 16'h9caa;
RsqrteLUT[6153] = 16'h9ca5;
RsqrteLUT[6154] = 16'h9ca1;
RsqrteLUT[6155] = 16'h9c9c;
RsqrteLUT[6156] = 16'h9c98;
RsqrteLUT[6157] = 16'h9c94;
RsqrteLUT[6158] = 16'h9c8f;
RsqrteLUT[6159] = 16'h9c8b;
RsqrteLUT[6160] = 16'h9c87;
RsqrteLUT[6161] = 16'h9c83;
RsqrteLUT[6162] = 16'h9c7f;
RsqrteLUT[6163] = 16'h9c7b;
RsqrteLUT[6164] = 16'h9c78;
RsqrteLUT[6165] = 16'h9c74;
RsqrteLUT[6166] = 16'h9c70;
RsqrteLUT[6167] = 16'h9c6d;
RsqrteLUT[6168] = 16'h9c69;
RsqrteLUT[6169] = 16'h9c66;
RsqrteLUT[6170] = 16'h9c62;
RsqrteLUT[6171] = 16'h9c5f;
RsqrteLUT[6172] = 16'h9c5b;
RsqrteLUT[6173] = 16'h9c58;
RsqrteLUT[6174] = 16'h9c55;
RsqrteLUT[6175] = 16'h9c52;
RsqrteLUT[6176] = 16'h9c4f;
RsqrteLUT[6177] = 16'h9c4c;
RsqrteLUT[6178] = 16'h9c49;
RsqrteLUT[6179] = 16'h9c46;
RsqrteLUT[6180] = 16'h9c43;
RsqrteLUT[6181] = 16'h9c40;
RsqrteLUT[6182] = 16'h9c3d;
RsqrteLUT[6183] = 16'h9c3a;
RsqrteLUT[6184] = 16'h9c38;
RsqrteLUT[6185] = 16'h9c35;
RsqrteLUT[6186] = 16'h9c32;
RsqrteLUT[6187] = 16'h9c2f;
RsqrteLUT[6188] = 16'h9c2d;
RsqrteLUT[6189] = 16'h9c2a;
RsqrteLUT[6190] = 16'h9c28;
RsqrteLUT[6191] = 16'h9c25;
RsqrteLUT[6192] = 16'h9c23;
RsqrteLUT[6193] = 16'h9c20;
RsqrteLUT[6194] = 16'h9c1e;
RsqrteLUT[6195] = 16'h9c1c;
RsqrteLUT[6196] = 16'h9c19;
RsqrteLUT[6197] = 16'h9c17;
RsqrteLUT[6198] = 16'h9c15;
RsqrteLUT[6199] = 16'h9c13;
RsqrteLUT[6200] = 16'h9c10;
RsqrteLUT[6201] = 16'h9c0e;
RsqrteLUT[6202] = 16'h9c0c;
RsqrteLUT[6203] = 16'h9c0a;
RsqrteLUT[6204] = 16'h9c08;
RsqrteLUT[6205] = 16'h9c06;
RsqrteLUT[6206] = 16'h9c04;
RsqrteLUT[6207] = 16'h9c02;
RsqrteLUT[6208] = 16'h9c00;
RsqrteLUT[6209] = 16'h9bf8;
RsqrteLUT[6210] = 16'h9bf0;
RsqrteLUT[6211] = 16'h9be8;
RsqrteLUT[6212] = 16'h9be1;
RsqrteLUT[6213] = 16'h9bda;
RsqrteLUT[6214] = 16'h9bd3;
RsqrteLUT[6215] = 16'h9bcc;
RsqrteLUT[6216] = 16'h9bc5;
RsqrteLUT[6217] = 16'h9bbe;
RsqrteLUT[6218] = 16'h9bb8;
RsqrteLUT[6219] = 16'h9bb1;
RsqrteLUT[6220] = 16'h9bab;
RsqrteLUT[6221] = 16'h9ba5;
RsqrteLUT[6222] = 16'h9b9f;
RsqrteLUT[6223] = 16'h9b99;
RsqrteLUT[6224] = 16'h9b93;
RsqrteLUT[6225] = 16'h9b8e;
RsqrteLUT[6226] = 16'h9b88;
RsqrteLUT[6227] = 16'h9b83;
RsqrteLUT[6228] = 16'h9b7d;
RsqrteLUT[6229] = 16'h9b78;
RsqrteLUT[6230] = 16'h9b73;
RsqrteLUT[6231] = 16'h9b6e;
RsqrteLUT[6232] = 16'h9b69;
RsqrteLUT[6233] = 16'h9b64;
RsqrteLUT[6234] = 16'h9b5f;
RsqrteLUT[6235] = 16'h9b5a;
RsqrteLUT[6236] = 16'h9b56;
RsqrteLUT[6237] = 16'h9b51;
RsqrteLUT[6238] = 16'h9b4c;
RsqrteLUT[6239] = 16'h9b48;
RsqrteLUT[6240] = 16'h9b44;
RsqrteLUT[6241] = 16'h9b3f;
RsqrteLUT[6242] = 16'h9b3b;
RsqrteLUT[6243] = 16'h9b37;
RsqrteLUT[6244] = 16'h9b33;
RsqrteLUT[6245] = 16'h9b2f;
RsqrteLUT[6246] = 16'h9b2b;
RsqrteLUT[6247] = 16'h9b27;
RsqrteLUT[6248] = 16'h9b23;
RsqrteLUT[6249] = 16'h9b1f;
RsqrteLUT[6250] = 16'h9b1b;
RsqrteLUT[6251] = 16'h9b17;
RsqrteLUT[6252] = 16'h9b14;
RsqrteLUT[6253] = 16'h9b10;
RsqrteLUT[6254] = 16'h9b0d;
RsqrteLUT[6255] = 16'h9b09;
RsqrteLUT[6256] = 16'h9b06;
RsqrteLUT[6257] = 16'h9b02;
RsqrteLUT[6258] = 16'h9aff;
RsqrteLUT[6259] = 16'h9afb;
RsqrteLUT[6260] = 16'h9af8;
RsqrteLUT[6261] = 16'h9af5;
RsqrteLUT[6262] = 16'h9af2;
RsqrteLUT[6263] = 16'h9aee;
RsqrteLUT[6264] = 16'h9aeb;
RsqrteLUT[6265] = 16'h9ae8;
RsqrteLUT[6266] = 16'h9ae5;
RsqrteLUT[6267] = 16'h9ae2;
RsqrteLUT[6268] = 16'h9adf;
RsqrteLUT[6269] = 16'h9adc;
RsqrteLUT[6270] = 16'h9ad9;
RsqrteLUT[6271] = 16'h9ad6;
RsqrteLUT[6272] = 16'h9ad4;
RsqrteLUT[6273] = 16'h9ace;
RsqrteLUT[6274] = 16'h9ac9;
RsqrteLUT[6275] = 16'h9ac3;
RsqrteLUT[6276] = 16'h9abe;
RsqrteLUT[6277] = 16'h9ab9;
RsqrteLUT[6278] = 16'h9ab4;
RsqrteLUT[6279] = 16'h9aaf;
RsqrteLUT[6280] = 16'h9aaa;
RsqrteLUT[6281] = 16'h9aa5;
RsqrteLUT[6282] = 16'h9aa1;
RsqrteLUT[6283] = 16'h9a9c;
RsqrteLUT[6284] = 16'h9a98;
RsqrteLUT[6285] = 16'h9a94;
RsqrteLUT[6286] = 16'h9a8f;
RsqrteLUT[6287] = 16'h9a8b;
RsqrteLUT[6288] = 16'h9a87;
RsqrteLUT[6289] = 16'h9a83;
RsqrteLUT[6290] = 16'h9a7f;
RsqrteLUT[6291] = 16'h9a7b;
RsqrteLUT[6292] = 16'h9a78;
RsqrteLUT[6293] = 16'h9a74;
RsqrteLUT[6294] = 16'h9a70;
RsqrteLUT[6295] = 16'h9a6d;
RsqrteLUT[6296] = 16'h9a69;
RsqrteLUT[6297] = 16'h9a66;
RsqrteLUT[6298] = 16'h9a62;
RsqrteLUT[6299] = 16'h9a5f;
RsqrteLUT[6300] = 16'h9a5b;
RsqrteLUT[6301] = 16'h9a58;
RsqrteLUT[6302] = 16'h9a55;
RsqrteLUT[6303] = 16'h9a52;
RsqrteLUT[6304] = 16'h9a4f;
RsqrteLUT[6305] = 16'h9a4c;
RsqrteLUT[6306] = 16'h9a49;
RsqrteLUT[6307] = 16'h9a46;
RsqrteLUT[6308] = 16'h9a43;
RsqrteLUT[6309] = 16'h9a40;
RsqrteLUT[6310] = 16'h9a3d;
RsqrteLUT[6311] = 16'h9a3a;
RsqrteLUT[6312] = 16'h9a38;
RsqrteLUT[6313] = 16'h9a35;
RsqrteLUT[6314] = 16'h9a32;
RsqrteLUT[6315] = 16'h9a2f;
RsqrteLUT[6316] = 16'h9a2d;
RsqrteLUT[6317] = 16'h9a2a;
RsqrteLUT[6318] = 16'h9a28;
RsqrteLUT[6319] = 16'h9a25;
RsqrteLUT[6320] = 16'h9a23;
RsqrteLUT[6321] = 16'h9a20;
RsqrteLUT[6322] = 16'h9a1e;
RsqrteLUT[6323] = 16'h9a1c;
RsqrteLUT[6324] = 16'h9a19;
RsqrteLUT[6325] = 16'h9a17;
RsqrteLUT[6326] = 16'h9a15;
RsqrteLUT[6327] = 16'h9a13;
RsqrteLUT[6328] = 16'h9a10;
RsqrteLUT[6329] = 16'h9a0e;
RsqrteLUT[6330] = 16'h9a0c;
RsqrteLUT[6331] = 16'h9a0a;
RsqrteLUT[6332] = 16'h9a08;
RsqrteLUT[6333] = 16'h9a06;
RsqrteLUT[6334] = 16'h9a04;
RsqrteLUT[6335] = 16'h9a02;
RsqrteLUT[6336] = 16'h9a00;
RsqrteLUT[6337] = 16'h99f8;
RsqrteLUT[6338] = 16'h99f0;
RsqrteLUT[6339] = 16'h99e8;
RsqrteLUT[6340] = 16'h99e1;
RsqrteLUT[6341] = 16'h99da;
RsqrteLUT[6342] = 16'h99d3;
RsqrteLUT[6343] = 16'h99cc;
RsqrteLUT[6344] = 16'h99c5;
RsqrteLUT[6345] = 16'h99be;
RsqrteLUT[6346] = 16'h99b8;
RsqrteLUT[6347] = 16'h99b1;
RsqrteLUT[6348] = 16'h99ab;
RsqrteLUT[6349] = 16'h99a5;
RsqrteLUT[6350] = 16'h999f;
RsqrteLUT[6351] = 16'h9999;
RsqrteLUT[6352] = 16'h9993;
RsqrteLUT[6353] = 16'h998e;
RsqrteLUT[6354] = 16'h9988;
RsqrteLUT[6355] = 16'h9983;
RsqrteLUT[6356] = 16'h997d;
RsqrteLUT[6357] = 16'h9978;
RsqrteLUT[6358] = 16'h9973;
RsqrteLUT[6359] = 16'h996e;
RsqrteLUT[6360] = 16'h9969;
RsqrteLUT[6361] = 16'h9964;
RsqrteLUT[6362] = 16'h995f;
RsqrteLUT[6363] = 16'h995a;
RsqrteLUT[6364] = 16'h9956;
RsqrteLUT[6365] = 16'h9951;
RsqrteLUT[6366] = 16'h994c;
RsqrteLUT[6367] = 16'h9948;
RsqrteLUT[6368] = 16'h9944;
RsqrteLUT[6369] = 16'h993f;
RsqrteLUT[6370] = 16'h993b;
RsqrteLUT[6371] = 16'h9937;
RsqrteLUT[6372] = 16'h9933;
RsqrteLUT[6373] = 16'h992f;
RsqrteLUT[6374] = 16'h992b;
RsqrteLUT[6375] = 16'h9927;
RsqrteLUT[6376] = 16'h9923;
RsqrteLUT[6377] = 16'h991f;
RsqrteLUT[6378] = 16'h991b;
RsqrteLUT[6379] = 16'h9917;
RsqrteLUT[6380] = 16'h9914;
RsqrteLUT[6381] = 16'h9910;
RsqrteLUT[6382] = 16'h990d;
RsqrteLUT[6383] = 16'h9909;
RsqrteLUT[6384] = 16'h9906;
RsqrteLUT[6385] = 16'h9902;
RsqrteLUT[6386] = 16'h98ff;
RsqrteLUT[6387] = 16'h98fb;
RsqrteLUT[6388] = 16'h98f8;
RsqrteLUT[6389] = 16'h98f5;
RsqrteLUT[6390] = 16'h98f2;
RsqrteLUT[6391] = 16'h98ee;
RsqrteLUT[6392] = 16'h98eb;
RsqrteLUT[6393] = 16'h98e8;
RsqrteLUT[6394] = 16'h98e5;
RsqrteLUT[6395] = 16'h98e2;
RsqrteLUT[6396] = 16'h98df;
RsqrteLUT[6397] = 16'h98dc;
RsqrteLUT[6398] = 16'h98d9;
RsqrteLUT[6399] = 16'h98d6;
RsqrteLUT[6400] = 16'h98d4;
RsqrteLUT[6401] = 16'h98ce;
RsqrteLUT[6402] = 16'h98c9;
RsqrteLUT[6403] = 16'h98c3;
RsqrteLUT[6404] = 16'h98be;
RsqrteLUT[6405] = 16'h98b9;
RsqrteLUT[6406] = 16'h98b4;
RsqrteLUT[6407] = 16'h98af;
RsqrteLUT[6408] = 16'h98aa;
RsqrteLUT[6409] = 16'h98a5;
RsqrteLUT[6410] = 16'h98a1;
RsqrteLUT[6411] = 16'h989c;
RsqrteLUT[6412] = 16'h9898;
RsqrteLUT[6413] = 16'h9894;
RsqrteLUT[6414] = 16'h988f;
RsqrteLUT[6415] = 16'h988b;
RsqrteLUT[6416] = 16'h9887;
RsqrteLUT[6417] = 16'h9883;
RsqrteLUT[6418] = 16'h987f;
RsqrteLUT[6419] = 16'h987b;
RsqrteLUT[6420] = 16'h9878;
RsqrteLUT[6421] = 16'h9874;
RsqrteLUT[6422] = 16'h9870;
RsqrteLUT[6423] = 16'h986d;
RsqrteLUT[6424] = 16'h9869;
RsqrteLUT[6425] = 16'h9866;
RsqrteLUT[6426] = 16'h9862;
RsqrteLUT[6427] = 16'h985f;
RsqrteLUT[6428] = 16'h985b;
RsqrteLUT[6429] = 16'h9858;
RsqrteLUT[6430] = 16'h9855;
RsqrteLUT[6431] = 16'h9852;
RsqrteLUT[6432] = 16'h984f;
RsqrteLUT[6433] = 16'h984c;
RsqrteLUT[6434] = 16'h9849;
RsqrteLUT[6435] = 16'h9846;
RsqrteLUT[6436] = 16'h9843;
RsqrteLUT[6437] = 16'h9840;
RsqrteLUT[6438] = 16'h983d;
RsqrteLUT[6439] = 16'h983a;
RsqrteLUT[6440] = 16'h9838;
RsqrteLUT[6441] = 16'h9835;
RsqrteLUT[6442] = 16'h9832;
RsqrteLUT[6443] = 16'h982f;
RsqrteLUT[6444] = 16'h982d;
RsqrteLUT[6445] = 16'h982a;
RsqrteLUT[6446] = 16'h9828;
RsqrteLUT[6447] = 16'h9825;
RsqrteLUT[6448] = 16'h9823;
RsqrteLUT[6449] = 16'h9820;
RsqrteLUT[6450] = 16'h981e;
RsqrteLUT[6451] = 16'h981c;
RsqrteLUT[6452] = 16'h9819;
RsqrteLUT[6453] = 16'h9817;
RsqrteLUT[6454] = 16'h9815;
RsqrteLUT[6455] = 16'h9813;
RsqrteLUT[6456] = 16'h9810;
RsqrteLUT[6457] = 16'h980e;
RsqrteLUT[6458] = 16'h980c;
RsqrteLUT[6459] = 16'h980a;
RsqrteLUT[6460] = 16'h9808;
RsqrteLUT[6461] = 16'h9806;
RsqrteLUT[6462] = 16'h9804;
RsqrteLUT[6463] = 16'h9802;
RsqrteLUT[6464] = 16'h9800;
RsqrteLUT[6465] = 16'h97f8;
RsqrteLUT[6466] = 16'h97f0;
RsqrteLUT[6467] = 16'h97e8;
RsqrteLUT[6468] = 16'h97e1;
RsqrteLUT[6469] = 16'h97da;
RsqrteLUT[6470] = 16'h97d3;
RsqrteLUT[6471] = 16'h97cc;
RsqrteLUT[6472] = 16'h97c5;
RsqrteLUT[6473] = 16'h97be;
RsqrteLUT[6474] = 16'h97b8;
RsqrteLUT[6475] = 16'h97b1;
RsqrteLUT[6476] = 16'h97ab;
RsqrteLUT[6477] = 16'h97a5;
RsqrteLUT[6478] = 16'h979f;
RsqrteLUT[6479] = 16'h9799;
RsqrteLUT[6480] = 16'h9793;
RsqrteLUT[6481] = 16'h978e;
RsqrteLUT[6482] = 16'h9788;
RsqrteLUT[6483] = 16'h9783;
RsqrteLUT[6484] = 16'h977d;
RsqrteLUT[6485] = 16'h9778;
RsqrteLUT[6486] = 16'h9773;
RsqrteLUT[6487] = 16'h976e;
RsqrteLUT[6488] = 16'h9769;
RsqrteLUT[6489] = 16'h9764;
RsqrteLUT[6490] = 16'h975f;
RsqrteLUT[6491] = 16'h975a;
RsqrteLUT[6492] = 16'h9756;
RsqrteLUT[6493] = 16'h9751;
RsqrteLUT[6494] = 16'h974c;
RsqrteLUT[6495] = 16'h9748;
RsqrteLUT[6496] = 16'h9744;
RsqrteLUT[6497] = 16'h973f;
RsqrteLUT[6498] = 16'h973b;
RsqrteLUT[6499] = 16'h9737;
RsqrteLUT[6500] = 16'h9733;
RsqrteLUT[6501] = 16'h972f;
RsqrteLUT[6502] = 16'h972b;
RsqrteLUT[6503] = 16'h9727;
RsqrteLUT[6504] = 16'h9723;
RsqrteLUT[6505] = 16'h971f;
RsqrteLUT[6506] = 16'h971b;
RsqrteLUT[6507] = 16'h9717;
RsqrteLUT[6508] = 16'h9714;
RsqrteLUT[6509] = 16'h9710;
RsqrteLUT[6510] = 16'h970d;
RsqrteLUT[6511] = 16'h9709;
RsqrteLUT[6512] = 16'h9706;
RsqrteLUT[6513] = 16'h9702;
RsqrteLUT[6514] = 16'h96ff;
RsqrteLUT[6515] = 16'h96fb;
RsqrteLUT[6516] = 16'h96f8;
RsqrteLUT[6517] = 16'h96f5;
RsqrteLUT[6518] = 16'h96f2;
RsqrteLUT[6519] = 16'h96ee;
RsqrteLUT[6520] = 16'h96eb;
RsqrteLUT[6521] = 16'h96e8;
RsqrteLUT[6522] = 16'h96e5;
RsqrteLUT[6523] = 16'h96e2;
RsqrteLUT[6524] = 16'h96df;
RsqrteLUT[6525] = 16'h96dc;
RsqrteLUT[6526] = 16'h96d9;
RsqrteLUT[6527] = 16'h96d6;
RsqrteLUT[6528] = 16'h96d4;
RsqrteLUT[6529] = 16'h96ce;
RsqrteLUT[6530] = 16'h96c9;
RsqrteLUT[6531] = 16'h96c3;
RsqrteLUT[6532] = 16'h96be;
RsqrteLUT[6533] = 16'h96b9;
RsqrteLUT[6534] = 16'h96b4;
RsqrteLUT[6535] = 16'h96af;
RsqrteLUT[6536] = 16'h96aa;
RsqrteLUT[6537] = 16'h96a5;
RsqrteLUT[6538] = 16'h96a1;
RsqrteLUT[6539] = 16'h969c;
RsqrteLUT[6540] = 16'h9698;
RsqrteLUT[6541] = 16'h9694;
RsqrteLUT[6542] = 16'h968f;
RsqrteLUT[6543] = 16'h968b;
RsqrteLUT[6544] = 16'h9687;
RsqrteLUT[6545] = 16'h9683;
RsqrteLUT[6546] = 16'h967f;
RsqrteLUT[6547] = 16'h967b;
RsqrteLUT[6548] = 16'h9678;
RsqrteLUT[6549] = 16'h9674;
RsqrteLUT[6550] = 16'h9670;
RsqrteLUT[6551] = 16'h966d;
RsqrteLUT[6552] = 16'h9669;
RsqrteLUT[6553] = 16'h9666;
RsqrteLUT[6554] = 16'h9662;
RsqrteLUT[6555] = 16'h965f;
RsqrteLUT[6556] = 16'h965b;
RsqrteLUT[6557] = 16'h9658;
RsqrteLUT[6558] = 16'h9655;
RsqrteLUT[6559] = 16'h9652;
RsqrteLUT[6560] = 16'h964f;
RsqrteLUT[6561] = 16'h964c;
RsqrteLUT[6562] = 16'h9649;
RsqrteLUT[6563] = 16'h9646;
RsqrteLUT[6564] = 16'h9643;
RsqrteLUT[6565] = 16'h9640;
RsqrteLUT[6566] = 16'h963d;
RsqrteLUT[6567] = 16'h963a;
RsqrteLUT[6568] = 16'h9638;
RsqrteLUT[6569] = 16'h9635;
RsqrteLUT[6570] = 16'h9632;
RsqrteLUT[6571] = 16'h962f;
RsqrteLUT[6572] = 16'h962d;
RsqrteLUT[6573] = 16'h962a;
RsqrteLUT[6574] = 16'h9628;
RsqrteLUT[6575] = 16'h9625;
RsqrteLUT[6576] = 16'h9623;
RsqrteLUT[6577] = 16'h9620;
RsqrteLUT[6578] = 16'h961e;
RsqrteLUT[6579] = 16'h961c;
RsqrteLUT[6580] = 16'h9619;
RsqrteLUT[6581] = 16'h9617;
RsqrteLUT[6582] = 16'h9615;
RsqrteLUT[6583] = 16'h9613;
RsqrteLUT[6584] = 16'h9610;
RsqrteLUT[6585] = 16'h960e;
RsqrteLUT[6586] = 16'h960c;
RsqrteLUT[6587] = 16'h960a;
RsqrteLUT[6588] = 16'h9608;
RsqrteLUT[6589] = 16'h9606;
RsqrteLUT[6590] = 16'h9604;
RsqrteLUT[6591] = 16'h9602;
RsqrteLUT[6592] = 16'h9600;
RsqrteLUT[6593] = 16'h95f8;
RsqrteLUT[6594] = 16'h95f0;
RsqrteLUT[6595] = 16'h95e8;
RsqrteLUT[6596] = 16'h95e1;
RsqrteLUT[6597] = 16'h95da;
RsqrteLUT[6598] = 16'h95d3;
RsqrteLUT[6599] = 16'h95cc;
RsqrteLUT[6600] = 16'h95c5;
RsqrteLUT[6601] = 16'h95be;
RsqrteLUT[6602] = 16'h95b8;
RsqrteLUT[6603] = 16'h95b1;
RsqrteLUT[6604] = 16'h95ab;
RsqrteLUT[6605] = 16'h95a5;
RsqrteLUT[6606] = 16'h959f;
RsqrteLUT[6607] = 16'h9599;
RsqrteLUT[6608] = 16'h9593;
RsqrteLUT[6609] = 16'h958e;
RsqrteLUT[6610] = 16'h9588;
RsqrteLUT[6611] = 16'h9583;
RsqrteLUT[6612] = 16'h957d;
RsqrteLUT[6613] = 16'h9578;
RsqrteLUT[6614] = 16'h9573;
RsqrteLUT[6615] = 16'h956e;
RsqrteLUT[6616] = 16'h9569;
RsqrteLUT[6617] = 16'h9564;
RsqrteLUT[6618] = 16'h955f;
RsqrteLUT[6619] = 16'h955a;
RsqrteLUT[6620] = 16'h9556;
RsqrteLUT[6621] = 16'h9551;
RsqrteLUT[6622] = 16'h954c;
RsqrteLUT[6623] = 16'h9548;
RsqrteLUT[6624] = 16'h9544;
RsqrteLUT[6625] = 16'h953f;
RsqrteLUT[6626] = 16'h953b;
RsqrteLUT[6627] = 16'h9537;
RsqrteLUT[6628] = 16'h9533;
RsqrteLUT[6629] = 16'h952f;
RsqrteLUT[6630] = 16'h952b;
RsqrteLUT[6631] = 16'h9527;
RsqrteLUT[6632] = 16'h9523;
RsqrteLUT[6633] = 16'h951f;
RsqrteLUT[6634] = 16'h951b;
RsqrteLUT[6635] = 16'h9517;
RsqrteLUT[6636] = 16'h9514;
RsqrteLUT[6637] = 16'h9510;
RsqrteLUT[6638] = 16'h950d;
RsqrteLUT[6639] = 16'h9509;
RsqrteLUT[6640] = 16'h9506;
RsqrteLUT[6641] = 16'h9502;
RsqrteLUT[6642] = 16'h94ff;
RsqrteLUT[6643] = 16'h94fb;
RsqrteLUT[6644] = 16'h94f8;
RsqrteLUT[6645] = 16'h94f5;
RsqrteLUT[6646] = 16'h94f2;
RsqrteLUT[6647] = 16'h94ee;
RsqrteLUT[6648] = 16'h94eb;
RsqrteLUT[6649] = 16'h94e8;
RsqrteLUT[6650] = 16'h94e5;
RsqrteLUT[6651] = 16'h94e2;
RsqrteLUT[6652] = 16'h94df;
RsqrteLUT[6653] = 16'h94dc;
RsqrteLUT[6654] = 16'h94d9;
RsqrteLUT[6655] = 16'h94d6;
RsqrteLUT[6656] = 16'h94d4;
RsqrteLUT[6657] = 16'h94ce;
RsqrteLUT[6658] = 16'h94c9;
RsqrteLUT[6659] = 16'h94c3;
RsqrteLUT[6660] = 16'h94be;
RsqrteLUT[6661] = 16'h94b9;
RsqrteLUT[6662] = 16'h94b4;
RsqrteLUT[6663] = 16'h94af;
RsqrteLUT[6664] = 16'h94aa;
RsqrteLUT[6665] = 16'h94a5;
RsqrteLUT[6666] = 16'h94a1;
RsqrteLUT[6667] = 16'h949c;
RsqrteLUT[6668] = 16'h9498;
RsqrteLUT[6669] = 16'h9494;
RsqrteLUT[6670] = 16'h948f;
RsqrteLUT[6671] = 16'h948b;
RsqrteLUT[6672] = 16'h9487;
RsqrteLUT[6673] = 16'h9483;
RsqrteLUT[6674] = 16'h947f;
RsqrteLUT[6675] = 16'h947b;
RsqrteLUT[6676] = 16'h9478;
RsqrteLUT[6677] = 16'h9474;
RsqrteLUT[6678] = 16'h9470;
RsqrteLUT[6679] = 16'h946d;
RsqrteLUT[6680] = 16'h9469;
RsqrteLUT[6681] = 16'h9466;
RsqrteLUT[6682] = 16'h9462;
RsqrteLUT[6683] = 16'h945f;
RsqrteLUT[6684] = 16'h945b;
RsqrteLUT[6685] = 16'h9458;
RsqrteLUT[6686] = 16'h9455;
RsqrteLUT[6687] = 16'h9452;
RsqrteLUT[6688] = 16'h944f;
RsqrteLUT[6689] = 16'h944c;
RsqrteLUT[6690] = 16'h9449;
RsqrteLUT[6691] = 16'h9446;
RsqrteLUT[6692] = 16'h9443;
RsqrteLUT[6693] = 16'h9440;
RsqrteLUT[6694] = 16'h943d;
RsqrteLUT[6695] = 16'h943a;
RsqrteLUT[6696] = 16'h9438;
RsqrteLUT[6697] = 16'h9435;
RsqrteLUT[6698] = 16'h9432;
RsqrteLUT[6699] = 16'h942f;
RsqrteLUT[6700] = 16'h942d;
RsqrteLUT[6701] = 16'h942a;
RsqrteLUT[6702] = 16'h9428;
RsqrteLUT[6703] = 16'h9425;
RsqrteLUT[6704] = 16'h9423;
RsqrteLUT[6705] = 16'h9420;
RsqrteLUT[6706] = 16'h941e;
RsqrteLUT[6707] = 16'h941c;
RsqrteLUT[6708] = 16'h9419;
RsqrteLUT[6709] = 16'h9417;
RsqrteLUT[6710] = 16'h9415;
RsqrteLUT[6711] = 16'h9413;
RsqrteLUT[6712] = 16'h9410;
RsqrteLUT[6713] = 16'h940e;
RsqrteLUT[6714] = 16'h940c;
RsqrteLUT[6715] = 16'h940a;
RsqrteLUT[6716] = 16'h9408;
RsqrteLUT[6717] = 16'h9406;
RsqrteLUT[6718] = 16'h9404;
RsqrteLUT[6719] = 16'h9402;
RsqrteLUT[6720] = 16'h9400;
RsqrteLUT[6721] = 16'h93f8;
RsqrteLUT[6722] = 16'h93f0;
RsqrteLUT[6723] = 16'h93e8;
RsqrteLUT[6724] = 16'h93e1;
RsqrteLUT[6725] = 16'h93da;
RsqrteLUT[6726] = 16'h93d3;
RsqrteLUT[6727] = 16'h93cc;
RsqrteLUT[6728] = 16'h93c5;
RsqrteLUT[6729] = 16'h93be;
RsqrteLUT[6730] = 16'h93b8;
RsqrteLUT[6731] = 16'h93b1;
RsqrteLUT[6732] = 16'h93ab;
RsqrteLUT[6733] = 16'h93a5;
RsqrteLUT[6734] = 16'h939f;
RsqrteLUT[6735] = 16'h9399;
RsqrteLUT[6736] = 16'h9393;
RsqrteLUT[6737] = 16'h938e;
RsqrteLUT[6738] = 16'h9388;
RsqrteLUT[6739] = 16'h9383;
RsqrteLUT[6740] = 16'h937d;
RsqrteLUT[6741] = 16'h9378;
RsqrteLUT[6742] = 16'h9373;
RsqrteLUT[6743] = 16'h936e;
RsqrteLUT[6744] = 16'h9369;
RsqrteLUT[6745] = 16'h9364;
RsqrteLUT[6746] = 16'h935f;
RsqrteLUT[6747] = 16'h935a;
RsqrteLUT[6748] = 16'h9356;
RsqrteLUT[6749] = 16'h9351;
RsqrteLUT[6750] = 16'h934c;
RsqrteLUT[6751] = 16'h9348;
RsqrteLUT[6752] = 16'h9344;
RsqrteLUT[6753] = 16'h933f;
RsqrteLUT[6754] = 16'h933b;
RsqrteLUT[6755] = 16'h9337;
RsqrteLUT[6756] = 16'h9333;
RsqrteLUT[6757] = 16'h932f;
RsqrteLUT[6758] = 16'h932b;
RsqrteLUT[6759] = 16'h9327;
RsqrteLUT[6760] = 16'h9323;
RsqrteLUT[6761] = 16'h931f;
RsqrteLUT[6762] = 16'h931b;
RsqrteLUT[6763] = 16'h9317;
RsqrteLUT[6764] = 16'h9314;
RsqrteLUT[6765] = 16'h9310;
RsqrteLUT[6766] = 16'h930d;
RsqrteLUT[6767] = 16'h9309;
RsqrteLUT[6768] = 16'h9306;
RsqrteLUT[6769] = 16'h9302;
RsqrteLUT[6770] = 16'h92ff;
RsqrteLUT[6771] = 16'h92fb;
RsqrteLUT[6772] = 16'h92f8;
RsqrteLUT[6773] = 16'h92f5;
RsqrteLUT[6774] = 16'h92f2;
RsqrteLUT[6775] = 16'h92ee;
RsqrteLUT[6776] = 16'h92eb;
RsqrteLUT[6777] = 16'h92e8;
RsqrteLUT[6778] = 16'h92e5;
RsqrteLUT[6779] = 16'h92e2;
RsqrteLUT[6780] = 16'h92df;
RsqrteLUT[6781] = 16'h92dc;
RsqrteLUT[6782] = 16'h92d9;
RsqrteLUT[6783] = 16'h92d6;
RsqrteLUT[6784] = 16'h92d4;
RsqrteLUT[6785] = 16'h92ce;
RsqrteLUT[6786] = 16'h92c9;
RsqrteLUT[6787] = 16'h92c3;
RsqrteLUT[6788] = 16'h92be;
RsqrteLUT[6789] = 16'h92b9;
RsqrteLUT[6790] = 16'h92b4;
RsqrteLUT[6791] = 16'h92af;
RsqrteLUT[6792] = 16'h92aa;
RsqrteLUT[6793] = 16'h92a5;
RsqrteLUT[6794] = 16'h92a1;
RsqrteLUT[6795] = 16'h929c;
RsqrteLUT[6796] = 16'h9298;
RsqrteLUT[6797] = 16'h9294;
RsqrteLUT[6798] = 16'h928f;
RsqrteLUT[6799] = 16'h928b;
RsqrteLUT[6800] = 16'h9287;
RsqrteLUT[6801] = 16'h9283;
RsqrteLUT[6802] = 16'h927f;
RsqrteLUT[6803] = 16'h927b;
RsqrteLUT[6804] = 16'h9278;
RsqrteLUT[6805] = 16'h9274;
RsqrteLUT[6806] = 16'h9270;
RsqrteLUT[6807] = 16'h926d;
RsqrteLUT[6808] = 16'h9269;
RsqrteLUT[6809] = 16'h9266;
RsqrteLUT[6810] = 16'h9262;
RsqrteLUT[6811] = 16'h925f;
RsqrteLUT[6812] = 16'h925b;
RsqrteLUT[6813] = 16'h9258;
RsqrteLUT[6814] = 16'h9255;
RsqrteLUT[6815] = 16'h9252;
RsqrteLUT[6816] = 16'h924f;
RsqrteLUT[6817] = 16'h924c;
RsqrteLUT[6818] = 16'h9249;
RsqrteLUT[6819] = 16'h9246;
RsqrteLUT[6820] = 16'h9243;
RsqrteLUT[6821] = 16'h9240;
RsqrteLUT[6822] = 16'h923d;
RsqrteLUT[6823] = 16'h923a;
RsqrteLUT[6824] = 16'h9238;
RsqrteLUT[6825] = 16'h9235;
RsqrteLUT[6826] = 16'h9232;
RsqrteLUT[6827] = 16'h922f;
RsqrteLUT[6828] = 16'h922d;
RsqrteLUT[6829] = 16'h922a;
RsqrteLUT[6830] = 16'h9228;
RsqrteLUT[6831] = 16'h9225;
RsqrteLUT[6832] = 16'h9223;
RsqrteLUT[6833] = 16'h9220;
RsqrteLUT[6834] = 16'h921e;
RsqrteLUT[6835] = 16'h921c;
RsqrteLUT[6836] = 16'h9219;
RsqrteLUT[6837] = 16'h9217;
RsqrteLUT[6838] = 16'h9215;
RsqrteLUT[6839] = 16'h9213;
RsqrteLUT[6840] = 16'h9210;
RsqrteLUT[6841] = 16'h920e;
RsqrteLUT[6842] = 16'h920c;
RsqrteLUT[6843] = 16'h920a;
RsqrteLUT[6844] = 16'h9208;
RsqrteLUT[6845] = 16'h9206;
RsqrteLUT[6846] = 16'h9204;
RsqrteLUT[6847] = 16'h9202;
RsqrteLUT[6848] = 16'h9200;
RsqrteLUT[6849] = 16'h91f8;
RsqrteLUT[6850] = 16'h91f0;
RsqrteLUT[6851] = 16'h91e8;
RsqrteLUT[6852] = 16'h91e1;
RsqrteLUT[6853] = 16'h91da;
RsqrteLUT[6854] = 16'h91d3;
RsqrteLUT[6855] = 16'h91cc;
RsqrteLUT[6856] = 16'h91c5;
RsqrteLUT[6857] = 16'h91be;
RsqrteLUT[6858] = 16'h91b8;
RsqrteLUT[6859] = 16'h91b1;
RsqrteLUT[6860] = 16'h91ab;
RsqrteLUT[6861] = 16'h91a5;
RsqrteLUT[6862] = 16'h919f;
RsqrteLUT[6863] = 16'h9199;
RsqrteLUT[6864] = 16'h9193;
RsqrteLUT[6865] = 16'h918e;
RsqrteLUT[6866] = 16'h9188;
RsqrteLUT[6867] = 16'h9183;
RsqrteLUT[6868] = 16'h917d;
RsqrteLUT[6869] = 16'h9178;
RsqrteLUT[6870] = 16'h9173;
RsqrteLUT[6871] = 16'h916e;
RsqrteLUT[6872] = 16'h9169;
RsqrteLUT[6873] = 16'h9164;
RsqrteLUT[6874] = 16'h915f;
RsqrteLUT[6875] = 16'h915a;
RsqrteLUT[6876] = 16'h9156;
RsqrteLUT[6877] = 16'h9151;
RsqrteLUT[6878] = 16'h914c;
RsqrteLUT[6879] = 16'h9148;
RsqrteLUT[6880] = 16'h9144;
RsqrteLUT[6881] = 16'h913f;
RsqrteLUT[6882] = 16'h913b;
RsqrteLUT[6883] = 16'h9137;
RsqrteLUT[6884] = 16'h9133;
RsqrteLUT[6885] = 16'h912f;
RsqrteLUT[6886] = 16'h912b;
RsqrteLUT[6887] = 16'h9127;
RsqrteLUT[6888] = 16'h9123;
RsqrteLUT[6889] = 16'h911f;
RsqrteLUT[6890] = 16'h911b;
RsqrteLUT[6891] = 16'h9117;
RsqrteLUT[6892] = 16'h9114;
RsqrteLUT[6893] = 16'h9110;
RsqrteLUT[6894] = 16'h910d;
RsqrteLUT[6895] = 16'h9109;
RsqrteLUT[6896] = 16'h9106;
RsqrteLUT[6897] = 16'h9102;
RsqrteLUT[6898] = 16'h90ff;
RsqrteLUT[6899] = 16'h90fb;
RsqrteLUT[6900] = 16'h90f8;
RsqrteLUT[6901] = 16'h90f5;
RsqrteLUT[6902] = 16'h90f2;
RsqrteLUT[6903] = 16'h90ee;
RsqrteLUT[6904] = 16'h90eb;
RsqrteLUT[6905] = 16'h90e8;
RsqrteLUT[6906] = 16'h90e5;
RsqrteLUT[6907] = 16'h90e2;
RsqrteLUT[6908] = 16'h90df;
RsqrteLUT[6909] = 16'h90dc;
RsqrteLUT[6910] = 16'h90d9;
RsqrteLUT[6911] = 16'h90d6;
RsqrteLUT[6912] = 16'h90d4;
RsqrteLUT[6913] = 16'h90ce;
RsqrteLUT[6914] = 16'h90c9;
RsqrteLUT[6915] = 16'h90c3;
RsqrteLUT[6916] = 16'h90be;
RsqrteLUT[6917] = 16'h90b9;
RsqrteLUT[6918] = 16'h90b4;
RsqrteLUT[6919] = 16'h90af;
RsqrteLUT[6920] = 16'h90aa;
RsqrteLUT[6921] = 16'h90a5;
RsqrteLUT[6922] = 16'h90a1;
RsqrteLUT[6923] = 16'h909c;
RsqrteLUT[6924] = 16'h9098;
RsqrteLUT[6925] = 16'h9094;
RsqrteLUT[6926] = 16'h908f;
RsqrteLUT[6927] = 16'h908b;
RsqrteLUT[6928] = 16'h9087;
RsqrteLUT[6929] = 16'h9083;
RsqrteLUT[6930] = 16'h907f;
RsqrteLUT[6931] = 16'h907b;
RsqrteLUT[6932] = 16'h9078;
RsqrteLUT[6933] = 16'h9074;
RsqrteLUT[6934] = 16'h9070;
RsqrteLUT[6935] = 16'h906d;
RsqrteLUT[6936] = 16'h9069;
RsqrteLUT[6937] = 16'h9066;
RsqrteLUT[6938] = 16'h9062;
RsqrteLUT[6939] = 16'h905f;
RsqrteLUT[6940] = 16'h905b;
RsqrteLUT[6941] = 16'h9058;
RsqrteLUT[6942] = 16'h9055;
RsqrteLUT[6943] = 16'h9052;
RsqrteLUT[6944] = 16'h904f;
RsqrteLUT[6945] = 16'h904c;
RsqrteLUT[6946] = 16'h9049;
RsqrteLUT[6947] = 16'h9046;
RsqrteLUT[6948] = 16'h9043;
RsqrteLUT[6949] = 16'h9040;
RsqrteLUT[6950] = 16'h903d;
RsqrteLUT[6951] = 16'h903a;
RsqrteLUT[6952] = 16'h9038;
RsqrteLUT[6953] = 16'h9035;
RsqrteLUT[6954] = 16'h9032;
RsqrteLUT[6955] = 16'h902f;
RsqrteLUT[6956] = 16'h902d;
RsqrteLUT[6957] = 16'h902a;
RsqrteLUT[6958] = 16'h9028;
RsqrteLUT[6959] = 16'h9025;
RsqrteLUT[6960] = 16'h9023;
RsqrteLUT[6961] = 16'h9020;
RsqrteLUT[6962] = 16'h901e;
RsqrteLUT[6963] = 16'h901c;
RsqrteLUT[6964] = 16'h9019;
RsqrteLUT[6965] = 16'h9017;
RsqrteLUT[6966] = 16'h9015;
RsqrteLUT[6967] = 16'h9013;
RsqrteLUT[6968] = 16'h9010;
RsqrteLUT[6969] = 16'h900e;
RsqrteLUT[6970] = 16'h900c;
RsqrteLUT[6971] = 16'h900a;
RsqrteLUT[6972] = 16'h9008;
RsqrteLUT[6973] = 16'h9006;
RsqrteLUT[6974] = 16'h9004;
RsqrteLUT[6975] = 16'h9002;
RsqrteLUT[6976] = 16'h9000;
RsqrteLUT[6977] = 16'h8ff8;
RsqrteLUT[6978] = 16'h8ff0;
RsqrteLUT[6979] = 16'h8fe8;
RsqrteLUT[6980] = 16'h8fe1;
RsqrteLUT[6981] = 16'h8fda;
RsqrteLUT[6982] = 16'h8fd3;
RsqrteLUT[6983] = 16'h8fcc;
RsqrteLUT[6984] = 16'h8fc5;
RsqrteLUT[6985] = 16'h8fbe;
RsqrteLUT[6986] = 16'h8fb8;
RsqrteLUT[6987] = 16'h8fb1;
RsqrteLUT[6988] = 16'h8fab;
RsqrteLUT[6989] = 16'h8fa5;
RsqrteLUT[6990] = 16'h8f9f;
RsqrteLUT[6991] = 16'h8f99;
RsqrteLUT[6992] = 16'h8f93;
RsqrteLUT[6993] = 16'h8f8e;
RsqrteLUT[6994] = 16'h8f88;
RsqrteLUT[6995] = 16'h8f83;
RsqrteLUT[6996] = 16'h8f7d;
RsqrteLUT[6997] = 16'h8f78;
RsqrteLUT[6998] = 16'h8f73;
RsqrteLUT[6999] = 16'h8f6e;
RsqrteLUT[7000] = 16'h8f69;
RsqrteLUT[7001] = 16'h8f64;
RsqrteLUT[7002] = 16'h8f5f;
RsqrteLUT[7003] = 16'h8f5a;
RsqrteLUT[7004] = 16'h8f56;
RsqrteLUT[7005] = 16'h8f51;
RsqrteLUT[7006] = 16'h8f4c;
RsqrteLUT[7007] = 16'h8f48;
RsqrteLUT[7008] = 16'h8f44;
RsqrteLUT[7009] = 16'h8f3f;
RsqrteLUT[7010] = 16'h8f3b;
RsqrteLUT[7011] = 16'h8f37;
RsqrteLUT[7012] = 16'h8f33;
RsqrteLUT[7013] = 16'h8f2f;
RsqrteLUT[7014] = 16'h8f2b;
RsqrteLUT[7015] = 16'h8f27;
RsqrteLUT[7016] = 16'h8f23;
RsqrteLUT[7017] = 16'h8f1f;
RsqrteLUT[7018] = 16'h8f1b;
RsqrteLUT[7019] = 16'h8f17;
RsqrteLUT[7020] = 16'h8f14;
RsqrteLUT[7021] = 16'h8f10;
RsqrteLUT[7022] = 16'h8f0d;
RsqrteLUT[7023] = 16'h8f09;
RsqrteLUT[7024] = 16'h8f06;
RsqrteLUT[7025] = 16'h8f02;
RsqrteLUT[7026] = 16'h8eff;
RsqrteLUT[7027] = 16'h8efb;
RsqrteLUT[7028] = 16'h8ef8;
RsqrteLUT[7029] = 16'h8ef5;
RsqrteLUT[7030] = 16'h8ef2;
RsqrteLUT[7031] = 16'h8eee;
RsqrteLUT[7032] = 16'h8eeb;
RsqrteLUT[7033] = 16'h8ee8;
RsqrteLUT[7034] = 16'h8ee5;
RsqrteLUT[7035] = 16'h8ee2;
RsqrteLUT[7036] = 16'h8edf;
RsqrteLUT[7037] = 16'h8edc;
RsqrteLUT[7038] = 16'h8ed9;
RsqrteLUT[7039] = 16'h8ed6;
RsqrteLUT[7040] = 16'h8ed4;
RsqrteLUT[7041] = 16'h8ece;
RsqrteLUT[7042] = 16'h8ec9;
RsqrteLUT[7043] = 16'h8ec3;
RsqrteLUT[7044] = 16'h8ebe;
RsqrteLUT[7045] = 16'h8eb9;
RsqrteLUT[7046] = 16'h8eb4;
RsqrteLUT[7047] = 16'h8eaf;
RsqrteLUT[7048] = 16'h8eaa;
RsqrteLUT[7049] = 16'h8ea5;
RsqrteLUT[7050] = 16'h8ea1;
RsqrteLUT[7051] = 16'h8e9c;
RsqrteLUT[7052] = 16'h8e98;
RsqrteLUT[7053] = 16'h8e94;
RsqrteLUT[7054] = 16'h8e8f;
RsqrteLUT[7055] = 16'h8e8b;
RsqrteLUT[7056] = 16'h8e87;
RsqrteLUT[7057] = 16'h8e83;
RsqrteLUT[7058] = 16'h8e7f;
RsqrteLUT[7059] = 16'h8e7b;
RsqrteLUT[7060] = 16'h8e78;
RsqrteLUT[7061] = 16'h8e74;
RsqrteLUT[7062] = 16'h8e70;
RsqrteLUT[7063] = 16'h8e6d;
RsqrteLUT[7064] = 16'h8e69;
RsqrteLUT[7065] = 16'h8e66;
RsqrteLUT[7066] = 16'h8e62;
RsqrteLUT[7067] = 16'h8e5f;
RsqrteLUT[7068] = 16'h8e5b;
RsqrteLUT[7069] = 16'h8e58;
RsqrteLUT[7070] = 16'h8e55;
RsqrteLUT[7071] = 16'h8e52;
RsqrteLUT[7072] = 16'h8e4f;
RsqrteLUT[7073] = 16'h8e4c;
RsqrteLUT[7074] = 16'h8e49;
RsqrteLUT[7075] = 16'h8e46;
RsqrteLUT[7076] = 16'h8e43;
RsqrteLUT[7077] = 16'h8e40;
RsqrteLUT[7078] = 16'h8e3d;
RsqrteLUT[7079] = 16'h8e3a;
RsqrteLUT[7080] = 16'h8e38;
RsqrteLUT[7081] = 16'h8e35;
RsqrteLUT[7082] = 16'h8e32;
RsqrteLUT[7083] = 16'h8e2f;
RsqrteLUT[7084] = 16'h8e2d;
RsqrteLUT[7085] = 16'h8e2a;
RsqrteLUT[7086] = 16'h8e28;
RsqrteLUT[7087] = 16'h8e25;
RsqrteLUT[7088] = 16'h8e23;
RsqrteLUT[7089] = 16'h8e20;
RsqrteLUT[7090] = 16'h8e1e;
RsqrteLUT[7091] = 16'h8e1c;
RsqrteLUT[7092] = 16'h8e19;
RsqrteLUT[7093] = 16'h8e17;
RsqrteLUT[7094] = 16'h8e15;
RsqrteLUT[7095] = 16'h8e13;
RsqrteLUT[7096] = 16'h8e10;
RsqrteLUT[7097] = 16'h8e0e;
RsqrteLUT[7098] = 16'h8e0c;
RsqrteLUT[7099] = 16'h8e0a;
RsqrteLUT[7100] = 16'h8e08;
RsqrteLUT[7101] = 16'h8e06;
RsqrteLUT[7102] = 16'h8e04;
RsqrteLUT[7103] = 16'h8e02;
RsqrteLUT[7104] = 16'h8e00;
RsqrteLUT[7105] = 16'h8df8;
RsqrteLUT[7106] = 16'h8df0;
RsqrteLUT[7107] = 16'h8de8;
RsqrteLUT[7108] = 16'h8de1;
RsqrteLUT[7109] = 16'h8dda;
RsqrteLUT[7110] = 16'h8dd3;
RsqrteLUT[7111] = 16'h8dcc;
RsqrteLUT[7112] = 16'h8dc5;
RsqrteLUT[7113] = 16'h8dbe;
RsqrteLUT[7114] = 16'h8db8;
RsqrteLUT[7115] = 16'h8db1;
RsqrteLUT[7116] = 16'h8dab;
RsqrteLUT[7117] = 16'h8da5;
RsqrteLUT[7118] = 16'h8d9f;
RsqrteLUT[7119] = 16'h8d99;
RsqrteLUT[7120] = 16'h8d93;
RsqrteLUT[7121] = 16'h8d8e;
RsqrteLUT[7122] = 16'h8d88;
RsqrteLUT[7123] = 16'h8d83;
RsqrteLUT[7124] = 16'h8d7d;
RsqrteLUT[7125] = 16'h8d78;
RsqrteLUT[7126] = 16'h8d73;
RsqrteLUT[7127] = 16'h8d6e;
RsqrteLUT[7128] = 16'h8d69;
RsqrteLUT[7129] = 16'h8d64;
RsqrteLUT[7130] = 16'h8d5f;
RsqrteLUT[7131] = 16'h8d5a;
RsqrteLUT[7132] = 16'h8d56;
RsqrteLUT[7133] = 16'h8d51;
RsqrteLUT[7134] = 16'h8d4c;
RsqrteLUT[7135] = 16'h8d48;
RsqrteLUT[7136] = 16'h8d44;
RsqrteLUT[7137] = 16'h8d3f;
RsqrteLUT[7138] = 16'h8d3b;
RsqrteLUT[7139] = 16'h8d37;
RsqrteLUT[7140] = 16'h8d33;
RsqrteLUT[7141] = 16'h8d2f;
RsqrteLUT[7142] = 16'h8d2b;
RsqrteLUT[7143] = 16'h8d27;
RsqrteLUT[7144] = 16'h8d23;
RsqrteLUT[7145] = 16'h8d1f;
RsqrteLUT[7146] = 16'h8d1b;
RsqrteLUT[7147] = 16'h8d17;
RsqrteLUT[7148] = 16'h8d14;
RsqrteLUT[7149] = 16'h8d10;
RsqrteLUT[7150] = 16'h8d0d;
RsqrteLUT[7151] = 16'h8d09;
RsqrteLUT[7152] = 16'h8d06;
RsqrteLUT[7153] = 16'h8d02;
RsqrteLUT[7154] = 16'h8cff;
RsqrteLUT[7155] = 16'h8cfb;
RsqrteLUT[7156] = 16'h8cf8;
RsqrteLUT[7157] = 16'h8cf5;
RsqrteLUT[7158] = 16'h8cf2;
RsqrteLUT[7159] = 16'h8cee;
RsqrteLUT[7160] = 16'h8ceb;
RsqrteLUT[7161] = 16'h8ce8;
RsqrteLUT[7162] = 16'h8ce5;
RsqrteLUT[7163] = 16'h8ce2;
RsqrteLUT[7164] = 16'h8cdf;
RsqrteLUT[7165] = 16'h8cdc;
RsqrteLUT[7166] = 16'h8cd9;
RsqrteLUT[7167] = 16'h8cd6;
RsqrteLUT[7168] = 16'h8cd4;
RsqrteLUT[7169] = 16'h8cce;
RsqrteLUT[7170] = 16'h8cc9;
RsqrteLUT[7171] = 16'h8cc3;
RsqrteLUT[7172] = 16'h8cbe;
RsqrteLUT[7173] = 16'h8cb9;
RsqrteLUT[7174] = 16'h8cb4;
RsqrteLUT[7175] = 16'h8caf;
RsqrteLUT[7176] = 16'h8caa;
RsqrteLUT[7177] = 16'h8ca5;
RsqrteLUT[7178] = 16'h8ca1;
RsqrteLUT[7179] = 16'h8c9c;
RsqrteLUT[7180] = 16'h8c98;
RsqrteLUT[7181] = 16'h8c94;
RsqrteLUT[7182] = 16'h8c8f;
RsqrteLUT[7183] = 16'h8c8b;
RsqrteLUT[7184] = 16'h8c87;
RsqrteLUT[7185] = 16'h8c83;
RsqrteLUT[7186] = 16'h8c7f;
RsqrteLUT[7187] = 16'h8c7b;
RsqrteLUT[7188] = 16'h8c78;
RsqrteLUT[7189] = 16'h8c74;
RsqrteLUT[7190] = 16'h8c70;
RsqrteLUT[7191] = 16'h8c6d;
RsqrteLUT[7192] = 16'h8c69;
RsqrteLUT[7193] = 16'h8c66;
RsqrteLUT[7194] = 16'h8c62;
RsqrteLUT[7195] = 16'h8c5f;
RsqrteLUT[7196] = 16'h8c5b;
RsqrteLUT[7197] = 16'h8c58;
RsqrteLUT[7198] = 16'h8c55;
RsqrteLUT[7199] = 16'h8c52;
RsqrteLUT[7200] = 16'h8c4f;
RsqrteLUT[7201] = 16'h8c4c;
RsqrteLUT[7202] = 16'h8c49;
RsqrteLUT[7203] = 16'h8c46;
RsqrteLUT[7204] = 16'h8c43;
RsqrteLUT[7205] = 16'h8c40;
RsqrteLUT[7206] = 16'h8c3d;
RsqrteLUT[7207] = 16'h8c3a;
RsqrteLUT[7208] = 16'h8c38;
RsqrteLUT[7209] = 16'h8c35;
RsqrteLUT[7210] = 16'h8c32;
RsqrteLUT[7211] = 16'h8c2f;
RsqrteLUT[7212] = 16'h8c2d;
RsqrteLUT[7213] = 16'h8c2a;
RsqrteLUT[7214] = 16'h8c28;
RsqrteLUT[7215] = 16'h8c25;
RsqrteLUT[7216] = 16'h8c23;
RsqrteLUT[7217] = 16'h8c20;
RsqrteLUT[7218] = 16'h8c1e;
RsqrteLUT[7219] = 16'h8c1c;
RsqrteLUT[7220] = 16'h8c19;
RsqrteLUT[7221] = 16'h8c17;
RsqrteLUT[7222] = 16'h8c15;
RsqrteLUT[7223] = 16'h8c13;
RsqrteLUT[7224] = 16'h8c10;
RsqrteLUT[7225] = 16'h8c0e;
RsqrteLUT[7226] = 16'h8c0c;
RsqrteLUT[7227] = 16'h8c0a;
RsqrteLUT[7228] = 16'h8c08;
RsqrteLUT[7229] = 16'h8c06;
RsqrteLUT[7230] = 16'h8c04;
RsqrteLUT[7231] = 16'h8c02;
RsqrteLUT[7232] = 16'h8c00;
RsqrteLUT[7233] = 16'h8bf8;
RsqrteLUT[7234] = 16'h8bf0;
RsqrteLUT[7235] = 16'h8be8;
RsqrteLUT[7236] = 16'h8be1;
RsqrteLUT[7237] = 16'h8bda;
RsqrteLUT[7238] = 16'h8bd3;
RsqrteLUT[7239] = 16'h8bcc;
RsqrteLUT[7240] = 16'h8bc5;
RsqrteLUT[7241] = 16'h8bbe;
RsqrteLUT[7242] = 16'h8bb8;
RsqrteLUT[7243] = 16'h8bb1;
RsqrteLUT[7244] = 16'h8bab;
RsqrteLUT[7245] = 16'h8ba5;
RsqrteLUT[7246] = 16'h8b9f;
RsqrteLUT[7247] = 16'h8b99;
RsqrteLUT[7248] = 16'h8b93;
RsqrteLUT[7249] = 16'h8b8e;
RsqrteLUT[7250] = 16'h8b88;
RsqrteLUT[7251] = 16'h8b83;
RsqrteLUT[7252] = 16'h8b7d;
RsqrteLUT[7253] = 16'h8b78;
RsqrteLUT[7254] = 16'h8b73;
RsqrteLUT[7255] = 16'h8b6e;
RsqrteLUT[7256] = 16'h8b69;
RsqrteLUT[7257] = 16'h8b64;
RsqrteLUT[7258] = 16'h8b5f;
RsqrteLUT[7259] = 16'h8b5a;
RsqrteLUT[7260] = 16'h8b56;
RsqrteLUT[7261] = 16'h8b51;
RsqrteLUT[7262] = 16'h8b4c;
RsqrteLUT[7263] = 16'h8b48;
RsqrteLUT[7264] = 16'h8b44;
RsqrteLUT[7265] = 16'h8b3f;
RsqrteLUT[7266] = 16'h8b3b;
RsqrteLUT[7267] = 16'h8b37;
RsqrteLUT[7268] = 16'h8b33;
RsqrteLUT[7269] = 16'h8b2f;
RsqrteLUT[7270] = 16'h8b2b;
RsqrteLUT[7271] = 16'h8b27;
RsqrteLUT[7272] = 16'h8b23;
RsqrteLUT[7273] = 16'h8b1f;
RsqrteLUT[7274] = 16'h8b1b;
RsqrteLUT[7275] = 16'h8b17;
RsqrteLUT[7276] = 16'h8b14;
RsqrteLUT[7277] = 16'h8b10;
RsqrteLUT[7278] = 16'h8b0d;
RsqrteLUT[7279] = 16'h8b09;
RsqrteLUT[7280] = 16'h8b06;
RsqrteLUT[7281] = 16'h8b02;
RsqrteLUT[7282] = 16'h8aff;
RsqrteLUT[7283] = 16'h8afb;
RsqrteLUT[7284] = 16'h8af8;
RsqrteLUT[7285] = 16'h8af5;
RsqrteLUT[7286] = 16'h8af2;
RsqrteLUT[7287] = 16'h8aee;
RsqrteLUT[7288] = 16'h8aeb;
RsqrteLUT[7289] = 16'h8ae8;
RsqrteLUT[7290] = 16'h8ae5;
RsqrteLUT[7291] = 16'h8ae2;
RsqrteLUT[7292] = 16'h8adf;
RsqrteLUT[7293] = 16'h8adc;
RsqrteLUT[7294] = 16'h8ad9;
RsqrteLUT[7295] = 16'h8ad6;
RsqrteLUT[7296] = 16'h8ad4;
RsqrteLUT[7297] = 16'h8ace;
RsqrteLUT[7298] = 16'h8ac9;
RsqrteLUT[7299] = 16'h8ac3;
RsqrteLUT[7300] = 16'h8abe;
RsqrteLUT[7301] = 16'h8ab9;
RsqrteLUT[7302] = 16'h8ab4;
RsqrteLUT[7303] = 16'h8aaf;
RsqrteLUT[7304] = 16'h8aaa;
RsqrteLUT[7305] = 16'h8aa5;
RsqrteLUT[7306] = 16'h8aa1;
RsqrteLUT[7307] = 16'h8a9c;
RsqrteLUT[7308] = 16'h8a98;
RsqrteLUT[7309] = 16'h8a94;
RsqrteLUT[7310] = 16'h8a8f;
RsqrteLUT[7311] = 16'h8a8b;
RsqrteLUT[7312] = 16'h8a87;
RsqrteLUT[7313] = 16'h8a83;
RsqrteLUT[7314] = 16'h8a7f;
RsqrteLUT[7315] = 16'h8a7b;
RsqrteLUT[7316] = 16'h8a78;
RsqrteLUT[7317] = 16'h8a74;
RsqrteLUT[7318] = 16'h8a70;
RsqrteLUT[7319] = 16'h8a6d;
RsqrteLUT[7320] = 16'h8a69;
RsqrteLUT[7321] = 16'h8a66;
RsqrteLUT[7322] = 16'h8a62;
RsqrteLUT[7323] = 16'h8a5f;
RsqrteLUT[7324] = 16'h8a5b;
RsqrteLUT[7325] = 16'h8a58;
RsqrteLUT[7326] = 16'h8a55;
RsqrteLUT[7327] = 16'h8a52;
RsqrteLUT[7328] = 16'h8a4f;
RsqrteLUT[7329] = 16'h8a4c;
RsqrteLUT[7330] = 16'h8a49;
RsqrteLUT[7331] = 16'h8a46;
RsqrteLUT[7332] = 16'h8a43;
RsqrteLUT[7333] = 16'h8a40;
RsqrteLUT[7334] = 16'h8a3d;
RsqrteLUT[7335] = 16'h8a3a;
RsqrteLUT[7336] = 16'h8a38;
RsqrteLUT[7337] = 16'h8a35;
RsqrteLUT[7338] = 16'h8a32;
RsqrteLUT[7339] = 16'h8a2f;
RsqrteLUT[7340] = 16'h8a2d;
RsqrteLUT[7341] = 16'h8a2a;
RsqrteLUT[7342] = 16'h8a28;
RsqrteLUT[7343] = 16'h8a25;
RsqrteLUT[7344] = 16'h8a23;
RsqrteLUT[7345] = 16'h8a20;
RsqrteLUT[7346] = 16'h8a1e;
RsqrteLUT[7347] = 16'h8a1c;
RsqrteLUT[7348] = 16'h8a19;
RsqrteLUT[7349] = 16'h8a17;
RsqrteLUT[7350] = 16'h8a15;
RsqrteLUT[7351] = 16'h8a13;
RsqrteLUT[7352] = 16'h8a10;
RsqrteLUT[7353] = 16'h8a0e;
RsqrteLUT[7354] = 16'h8a0c;
RsqrteLUT[7355] = 16'h8a0a;
RsqrteLUT[7356] = 16'h8a08;
RsqrteLUT[7357] = 16'h8a06;
RsqrteLUT[7358] = 16'h8a04;
RsqrteLUT[7359] = 16'h8a02;
RsqrteLUT[7360] = 16'h8a00;
RsqrteLUT[7361] = 16'h89f8;
RsqrteLUT[7362] = 16'h89f0;
RsqrteLUT[7363] = 16'h89e8;
RsqrteLUT[7364] = 16'h89e1;
RsqrteLUT[7365] = 16'h89da;
RsqrteLUT[7366] = 16'h89d3;
RsqrteLUT[7367] = 16'h89cc;
RsqrteLUT[7368] = 16'h89c5;
RsqrteLUT[7369] = 16'h89be;
RsqrteLUT[7370] = 16'h89b8;
RsqrteLUT[7371] = 16'h89b1;
RsqrteLUT[7372] = 16'h89ab;
RsqrteLUT[7373] = 16'h89a5;
RsqrteLUT[7374] = 16'h899f;
RsqrteLUT[7375] = 16'h8999;
RsqrteLUT[7376] = 16'h8993;
RsqrteLUT[7377] = 16'h898e;
RsqrteLUT[7378] = 16'h8988;
RsqrteLUT[7379] = 16'h8983;
RsqrteLUT[7380] = 16'h897d;
RsqrteLUT[7381] = 16'h8978;
RsqrteLUT[7382] = 16'h8973;
RsqrteLUT[7383] = 16'h896e;
RsqrteLUT[7384] = 16'h8969;
RsqrteLUT[7385] = 16'h8964;
RsqrteLUT[7386] = 16'h895f;
RsqrteLUT[7387] = 16'h895a;
RsqrteLUT[7388] = 16'h8956;
RsqrteLUT[7389] = 16'h8951;
RsqrteLUT[7390] = 16'h894c;
RsqrteLUT[7391] = 16'h8948;
RsqrteLUT[7392] = 16'h8944;
RsqrteLUT[7393] = 16'h893f;
RsqrteLUT[7394] = 16'h893b;
RsqrteLUT[7395] = 16'h8937;
RsqrteLUT[7396] = 16'h8933;
RsqrteLUT[7397] = 16'h892f;
RsqrteLUT[7398] = 16'h892b;
RsqrteLUT[7399] = 16'h8927;
RsqrteLUT[7400] = 16'h8923;
RsqrteLUT[7401] = 16'h891f;
RsqrteLUT[7402] = 16'h891b;
RsqrteLUT[7403] = 16'h8917;
RsqrteLUT[7404] = 16'h8914;
RsqrteLUT[7405] = 16'h8910;
RsqrteLUT[7406] = 16'h890d;
RsqrteLUT[7407] = 16'h8909;
RsqrteLUT[7408] = 16'h8906;
RsqrteLUT[7409] = 16'h8902;
RsqrteLUT[7410] = 16'h88ff;
RsqrteLUT[7411] = 16'h88fb;
RsqrteLUT[7412] = 16'h88f8;
RsqrteLUT[7413] = 16'h88f5;
RsqrteLUT[7414] = 16'h88f2;
RsqrteLUT[7415] = 16'h88ee;
RsqrteLUT[7416] = 16'h88eb;
RsqrteLUT[7417] = 16'h88e8;
RsqrteLUT[7418] = 16'h88e5;
RsqrteLUT[7419] = 16'h88e2;
RsqrteLUT[7420] = 16'h88df;
RsqrteLUT[7421] = 16'h88dc;
RsqrteLUT[7422] = 16'h88d9;
RsqrteLUT[7423] = 16'h88d6;
RsqrteLUT[7424] = 16'h88d4;
RsqrteLUT[7425] = 16'h88ce;
RsqrteLUT[7426] = 16'h88c9;
RsqrteLUT[7427] = 16'h88c3;
RsqrteLUT[7428] = 16'h88be;
RsqrteLUT[7429] = 16'h88b9;
RsqrteLUT[7430] = 16'h88b4;
RsqrteLUT[7431] = 16'h88af;
RsqrteLUT[7432] = 16'h88aa;
RsqrteLUT[7433] = 16'h88a5;
RsqrteLUT[7434] = 16'h88a1;
RsqrteLUT[7435] = 16'h889c;
RsqrteLUT[7436] = 16'h8898;
RsqrteLUT[7437] = 16'h8894;
RsqrteLUT[7438] = 16'h888f;
RsqrteLUT[7439] = 16'h888b;
RsqrteLUT[7440] = 16'h8887;
RsqrteLUT[7441] = 16'h8883;
RsqrteLUT[7442] = 16'h887f;
RsqrteLUT[7443] = 16'h887b;
RsqrteLUT[7444] = 16'h8878;
RsqrteLUT[7445] = 16'h8874;
RsqrteLUT[7446] = 16'h8870;
RsqrteLUT[7447] = 16'h886d;
RsqrteLUT[7448] = 16'h8869;
RsqrteLUT[7449] = 16'h8866;
RsqrteLUT[7450] = 16'h8862;
RsqrteLUT[7451] = 16'h885f;
RsqrteLUT[7452] = 16'h885b;
RsqrteLUT[7453] = 16'h8858;
RsqrteLUT[7454] = 16'h8855;
RsqrteLUT[7455] = 16'h8852;
RsqrteLUT[7456] = 16'h884f;
RsqrteLUT[7457] = 16'h884c;
RsqrteLUT[7458] = 16'h8849;
RsqrteLUT[7459] = 16'h8846;
RsqrteLUT[7460] = 16'h8843;
RsqrteLUT[7461] = 16'h8840;
RsqrteLUT[7462] = 16'h883d;
RsqrteLUT[7463] = 16'h883a;
RsqrteLUT[7464] = 16'h8838;
RsqrteLUT[7465] = 16'h8835;
RsqrteLUT[7466] = 16'h8832;
RsqrteLUT[7467] = 16'h882f;
RsqrteLUT[7468] = 16'h882d;
RsqrteLUT[7469] = 16'h882a;
RsqrteLUT[7470] = 16'h8828;
RsqrteLUT[7471] = 16'h8825;
RsqrteLUT[7472] = 16'h8823;
RsqrteLUT[7473] = 16'h8820;
RsqrteLUT[7474] = 16'h881e;
RsqrteLUT[7475] = 16'h881c;
RsqrteLUT[7476] = 16'h8819;
RsqrteLUT[7477] = 16'h8817;
RsqrteLUT[7478] = 16'h8815;
RsqrteLUT[7479] = 16'h8813;
RsqrteLUT[7480] = 16'h8810;
RsqrteLUT[7481] = 16'h880e;
RsqrteLUT[7482] = 16'h880c;
RsqrteLUT[7483] = 16'h880a;
RsqrteLUT[7484] = 16'h8808;
RsqrteLUT[7485] = 16'h8806;
RsqrteLUT[7486] = 16'h8804;
RsqrteLUT[7487] = 16'h8802;
RsqrteLUT[7488] = 16'h8800;
RsqrteLUT[7489] = 16'h87f8;
RsqrteLUT[7490] = 16'h87f0;
RsqrteLUT[7491] = 16'h87e8;
RsqrteLUT[7492] = 16'h87e1;
RsqrteLUT[7493] = 16'h87da;
RsqrteLUT[7494] = 16'h87d3;
RsqrteLUT[7495] = 16'h87cc;
RsqrteLUT[7496] = 16'h87c5;
RsqrteLUT[7497] = 16'h87be;
RsqrteLUT[7498] = 16'h87b8;
RsqrteLUT[7499] = 16'h87b1;
RsqrteLUT[7500] = 16'h87ab;
RsqrteLUT[7501] = 16'h87a5;
RsqrteLUT[7502] = 16'h879f;
RsqrteLUT[7503] = 16'h8799;
RsqrteLUT[7504] = 16'h8793;
RsqrteLUT[7505] = 16'h878e;
RsqrteLUT[7506] = 16'h8788;
RsqrteLUT[7507] = 16'h8783;
RsqrteLUT[7508] = 16'h877d;
RsqrteLUT[7509] = 16'h8778;
RsqrteLUT[7510] = 16'h8773;
RsqrteLUT[7511] = 16'h876e;
RsqrteLUT[7512] = 16'h8769;
RsqrteLUT[7513] = 16'h8764;
RsqrteLUT[7514] = 16'h875f;
RsqrteLUT[7515] = 16'h875a;
RsqrteLUT[7516] = 16'h8756;
RsqrteLUT[7517] = 16'h8751;
RsqrteLUT[7518] = 16'h874c;
RsqrteLUT[7519] = 16'h8748;
RsqrteLUT[7520] = 16'h8744;
RsqrteLUT[7521] = 16'h873f;
RsqrteLUT[7522] = 16'h873b;
RsqrteLUT[7523] = 16'h8737;
RsqrteLUT[7524] = 16'h8733;
RsqrteLUT[7525] = 16'h872f;
RsqrteLUT[7526] = 16'h872b;
RsqrteLUT[7527] = 16'h8727;
RsqrteLUT[7528] = 16'h8723;
RsqrteLUT[7529] = 16'h871f;
RsqrteLUT[7530] = 16'h871b;
RsqrteLUT[7531] = 16'h8717;
RsqrteLUT[7532] = 16'h8714;
RsqrteLUT[7533] = 16'h8710;
RsqrteLUT[7534] = 16'h870d;
RsqrteLUT[7535] = 16'h8709;
RsqrteLUT[7536] = 16'h8706;
RsqrteLUT[7537] = 16'h8702;
RsqrteLUT[7538] = 16'h86ff;
RsqrteLUT[7539] = 16'h86fb;
RsqrteLUT[7540] = 16'h86f8;
RsqrteLUT[7541] = 16'h86f5;
RsqrteLUT[7542] = 16'h86f2;
RsqrteLUT[7543] = 16'h86ee;
RsqrteLUT[7544] = 16'h86eb;
RsqrteLUT[7545] = 16'h86e8;
RsqrteLUT[7546] = 16'h86e5;
RsqrteLUT[7547] = 16'h86e2;
RsqrteLUT[7548] = 16'h86df;
RsqrteLUT[7549] = 16'h86dc;
RsqrteLUT[7550] = 16'h86d9;
RsqrteLUT[7551] = 16'h86d6;
RsqrteLUT[7552] = 16'h86d4;
RsqrteLUT[7553] = 16'h86ce;
RsqrteLUT[7554] = 16'h86c9;
RsqrteLUT[7555] = 16'h86c3;
RsqrteLUT[7556] = 16'h86be;
RsqrteLUT[7557] = 16'h86b9;
RsqrteLUT[7558] = 16'h86b4;
RsqrteLUT[7559] = 16'h86af;
RsqrteLUT[7560] = 16'h86aa;
RsqrteLUT[7561] = 16'h86a5;
RsqrteLUT[7562] = 16'h86a1;
RsqrteLUT[7563] = 16'h869c;
RsqrteLUT[7564] = 16'h8698;
RsqrteLUT[7565] = 16'h8694;
RsqrteLUT[7566] = 16'h868f;
RsqrteLUT[7567] = 16'h868b;
RsqrteLUT[7568] = 16'h8687;
RsqrteLUT[7569] = 16'h8683;
RsqrteLUT[7570] = 16'h867f;
RsqrteLUT[7571] = 16'h867b;
RsqrteLUT[7572] = 16'h8678;
RsqrteLUT[7573] = 16'h8674;
RsqrteLUT[7574] = 16'h8670;
RsqrteLUT[7575] = 16'h866d;
RsqrteLUT[7576] = 16'h8669;
RsqrteLUT[7577] = 16'h8666;
RsqrteLUT[7578] = 16'h8662;
RsqrteLUT[7579] = 16'h865f;
RsqrteLUT[7580] = 16'h865b;
RsqrteLUT[7581] = 16'h8658;
RsqrteLUT[7582] = 16'h8655;
RsqrteLUT[7583] = 16'h8652;
RsqrteLUT[7584] = 16'h864f;
RsqrteLUT[7585] = 16'h864c;
RsqrteLUT[7586] = 16'h8649;
RsqrteLUT[7587] = 16'h8646;
RsqrteLUT[7588] = 16'h8643;
RsqrteLUT[7589] = 16'h8640;
RsqrteLUT[7590] = 16'h863d;
RsqrteLUT[7591] = 16'h863a;
RsqrteLUT[7592] = 16'h8638;
RsqrteLUT[7593] = 16'h8635;
RsqrteLUT[7594] = 16'h8632;
RsqrteLUT[7595] = 16'h862f;
RsqrteLUT[7596] = 16'h862d;
RsqrteLUT[7597] = 16'h862a;
RsqrteLUT[7598] = 16'h8628;
RsqrteLUT[7599] = 16'h8625;
RsqrteLUT[7600] = 16'h8623;
RsqrteLUT[7601] = 16'h8620;
RsqrteLUT[7602] = 16'h861e;
RsqrteLUT[7603] = 16'h861c;
RsqrteLUT[7604] = 16'h8619;
RsqrteLUT[7605] = 16'h8617;
RsqrteLUT[7606] = 16'h8615;
RsqrteLUT[7607] = 16'h8613;
RsqrteLUT[7608] = 16'h8610;
RsqrteLUT[7609] = 16'h860e;
RsqrteLUT[7610] = 16'h860c;
RsqrteLUT[7611] = 16'h860a;
RsqrteLUT[7612] = 16'h8608;
RsqrteLUT[7613] = 16'h8606;
RsqrteLUT[7614] = 16'h8604;
RsqrteLUT[7615] = 16'h8602;
RsqrteLUT[7616] = 16'h8600;
RsqrteLUT[7617] = 16'h85f8;
RsqrteLUT[7618] = 16'h85f0;
RsqrteLUT[7619] = 16'h85e8;
RsqrteLUT[7620] = 16'h85e1;
RsqrteLUT[7621] = 16'h85da;
RsqrteLUT[7622] = 16'h85d3;
RsqrteLUT[7623] = 16'h85cc;
RsqrteLUT[7624] = 16'h85c5;
RsqrteLUT[7625] = 16'h85be;
RsqrteLUT[7626] = 16'h85b8;
RsqrteLUT[7627] = 16'h85b1;
RsqrteLUT[7628] = 16'h85ab;
RsqrteLUT[7629] = 16'h85a5;
RsqrteLUT[7630] = 16'h859f;
RsqrteLUT[7631] = 16'h8599;
RsqrteLUT[7632] = 16'h8593;
RsqrteLUT[7633] = 16'h858e;
RsqrteLUT[7634] = 16'h8588;
RsqrteLUT[7635] = 16'h8583;
RsqrteLUT[7636] = 16'h857d;
RsqrteLUT[7637] = 16'h8578;
RsqrteLUT[7638] = 16'h8573;
RsqrteLUT[7639] = 16'h856e;
RsqrteLUT[7640] = 16'h8569;
RsqrteLUT[7641] = 16'h8564;
RsqrteLUT[7642] = 16'h855f;
RsqrteLUT[7643] = 16'h855a;
RsqrteLUT[7644] = 16'h8556;
RsqrteLUT[7645] = 16'h8551;
RsqrteLUT[7646] = 16'h854c;
RsqrteLUT[7647] = 16'h8548;
RsqrteLUT[7648] = 16'h8544;
RsqrteLUT[7649] = 16'h853f;
RsqrteLUT[7650] = 16'h853b;
RsqrteLUT[7651] = 16'h8537;
RsqrteLUT[7652] = 16'h8533;
RsqrteLUT[7653] = 16'h852f;
RsqrteLUT[7654] = 16'h852b;
RsqrteLUT[7655] = 16'h8527;
RsqrteLUT[7656] = 16'h8523;
RsqrteLUT[7657] = 16'h851f;
RsqrteLUT[7658] = 16'h851b;
RsqrteLUT[7659] = 16'h8517;
RsqrteLUT[7660] = 16'h8514;
RsqrteLUT[7661] = 16'h8510;
RsqrteLUT[7662] = 16'h850d;
RsqrteLUT[7663] = 16'h8509;
RsqrteLUT[7664] = 16'h8506;
RsqrteLUT[7665] = 16'h8502;
RsqrteLUT[7666] = 16'h84ff;
RsqrteLUT[7667] = 16'h84fb;
RsqrteLUT[7668] = 16'h84f8;
RsqrteLUT[7669] = 16'h84f5;
RsqrteLUT[7670] = 16'h84f2;
RsqrteLUT[7671] = 16'h84ee;
RsqrteLUT[7672] = 16'h84eb;
RsqrteLUT[7673] = 16'h84e8;
RsqrteLUT[7674] = 16'h84e5;
RsqrteLUT[7675] = 16'h84e2;
RsqrteLUT[7676] = 16'h84df;
RsqrteLUT[7677] = 16'h84dc;
RsqrteLUT[7678] = 16'h84d9;
RsqrteLUT[7679] = 16'h84d6;
RsqrteLUT[7680] = 16'h84d4;
RsqrteLUT[7681] = 16'h84ce;
RsqrteLUT[7682] = 16'h84c9;
RsqrteLUT[7683] = 16'h84c3;
RsqrteLUT[7684] = 16'h84be;
RsqrteLUT[7685] = 16'h84b9;
RsqrteLUT[7686] = 16'h84b4;
RsqrteLUT[7687] = 16'h84af;
RsqrteLUT[7688] = 16'h84aa;
RsqrteLUT[7689] = 16'h84a5;
RsqrteLUT[7690] = 16'h84a1;
RsqrteLUT[7691] = 16'h849c;
RsqrteLUT[7692] = 16'h8498;
RsqrteLUT[7693] = 16'h8494;
RsqrteLUT[7694] = 16'h848f;
RsqrteLUT[7695] = 16'h848b;
RsqrteLUT[7696] = 16'h8487;
RsqrteLUT[7697] = 16'h8483;
RsqrteLUT[7698] = 16'h847f;
RsqrteLUT[7699] = 16'h847b;
RsqrteLUT[7700] = 16'h8478;
RsqrteLUT[7701] = 16'h8474;
RsqrteLUT[7702] = 16'h8470;
RsqrteLUT[7703] = 16'h846d;
RsqrteLUT[7704] = 16'h8469;
RsqrteLUT[7705] = 16'h8466;
RsqrteLUT[7706] = 16'h8462;
RsqrteLUT[7707] = 16'h845f;
RsqrteLUT[7708] = 16'h845b;
RsqrteLUT[7709] = 16'h8458;
RsqrteLUT[7710] = 16'h8455;
RsqrteLUT[7711] = 16'h8452;
RsqrteLUT[7712] = 16'h844f;
RsqrteLUT[7713] = 16'h844c;
RsqrteLUT[7714] = 16'h8449;
RsqrteLUT[7715] = 16'h8446;
RsqrteLUT[7716] = 16'h8443;
RsqrteLUT[7717] = 16'h8440;
RsqrteLUT[7718] = 16'h843d;
RsqrteLUT[7719] = 16'h843a;
RsqrteLUT[7720] = 16'h8438;
RsqrteLUT[7721] = 16'h8435;
RsqrteLUT[7722] = 16'h8432;
RsqrteLUT[7723] = 16'h842f;
RsqrteLUT[7724] = 16'h842d;
RsqrteLUT[7725] = 16'h842a;
RsqrteLUT[7726] = 16'h8428;
RsqrteLUT[7727] = 16'h8425;
RsqrteLUT[7728] = 16'h8423;
RsqrteLUT[7729] = 16'h8420;
RsqrteLUT[7730] = 16'h841e;
RsqrteLUT[7731] = 16'h841c;
RsqrteLUT[7732] = 16'h8419;
RsqrteLUT[7733] = 16'h8417;
RsqrteLUT[7734] = 16'h8415;
RsqrteLUT[7735] = 16'h8413;
RsqrteLUT[7736] = 16'h8410;
RsqrteLUT[7737] = 16'h840e;
RsqrteLUT[7738] = 16'h840c;
RsqrteLUT[7739] = 16'h840a;
RsqrteLUT[7740] = 16'h8408;
RsqrteLUT[7741] = 16'h8406;
RsqrteLUT[7742] = 16'h8404;
RsqrteLUT[7743] = 16'h8402;
RsqrteLUT[7744] = 16'h8400;
RsqrteLUT[7745] = 16'h83f8;
RsqrteLUT[7746] = 16'h83f0;
RsqrteLUT[7747] = 16'h83e8;
RsqrteLUT[7748] = 16'h83e1;
RsqrteLUT[7749] = 16'h83da;
RsqrteLUT[7750] = 16'h83d3;
RsqrteLUT[7751] = 16'h83cc;
RsqrteLUT[7752] = 16'h83c5;
RsqrteLUT[7753] = 16'h83be;
RsqrteLUT[7754] = 16'h83b8;
RsqrteLUT[7755] = 16'h83b1;
RsqrteLUT[7756] = 16'h83ab;
RsqrteLUT[7757] = 16'h83a5;
RsqrteLUT[7758] = 16'h839f;
RsqrteLUT[7759] = 16'h8399;
RsqrteLUT[7760] = 16'h8393;
RsqrteLUT[7761] = 16'h838e;
RsqrteLUT[7762] = 16'h8388;
RsqrteLUT[7763] = 16'h8383;
RsqrteLUT[7764] = 16'h837d;
RsqrteLUT[7765] = 16'h8378;
RsqrteLUT[7766] = 16'h8373;
RsqrteLUT[7767] = 16'h836e;
RsqrteLUT[7768] = 16'h8369;
RsqrteLUT[7769] = 16'h8364;
RsqrteLUT[7770] = 16'h835f;
RsqrteLUT[7771] = 16'h835a;
RsqrteLUT[7772] = 16'h8356;
RsqrteLUT[7773] = 16'h8351;
RsqrteLUT[7774] = 16'h834c;
RsqrteLUT[7775] = 16'h8348;
RsqrteLUT[7776] = 16'h8344;
RsqrteLUT[7777] = 16'h833f;
RsqrteLUT[7778] = 16'h833b;
RsqrteLUT[7779] = 16'h8337;
RsqrteLUT[7780] = 16'h8333;
RsqrteLUT[7781] = 16'h832f;
RsqrteLUT[7782] = 16'h832b;
RsqrteLUT[7783] = 16'h8327;
RsqrteLUT[7784] = 16'h8323;
RsqrteLUT[7785] = 16'h831f;
RsqrteLUT[7786] = 16'h831b;
RsqrteLUT[7787] = 16'h8317;
RsqrteLUT[7788] = 16'h8314;
RsqrteLUT[7789] = 16'h8310;
RsqrteLUT[7790] = 16'h830d;
RsqrteLUT[7791] = 16'h8309;
RsqrteLUT[7792] = 16'h8306;
RsqrteLUT[7793] = 16'h8302;
RsqrteLUT[7794] = 16'h82ff;
RsqrteLUT[7795] = 16'h82fb;
RsqrteLUT[7796] = 16'h82f8;
RsqrteLUT[7797] = 16'h82f5;
RsqrteLUT[7798] = 16'h82f2;
RsqrteLUT[7799] = 16'h82ee;
RsqrteLUT[7800] = 16'h82eb;
RsqrteLUT[7801] = 16'h82e8;
RsqrteLUT[7802] = 16'h82e5;
RsqrteLUT[7803] = 16'h82e2;
RsqrteLUT[7804] = 16'h82df;
RsqrteLUT[7805] = 16'h82dc;
RsqrteLUT[7806] = 16'h82d9;
RsqrteLUT[7807] = 16'h82d6;
RsqrteLUT[7808] = 16'h82d4;
RsqrteLUT[7809] = 16'h82ce;
RsqrteLUT[7810] = 16'h82c9;
RsqrteLUT[7811] = 16'h82c3;
RsqrteLUT[7812] = 16'h82be;
RsqrteLUT[7813] = 16'h82b9;
RsqrteLUT[7814] = 16'h82b4;
RsqrteLUT[7815] = 16'h82af;
RsqrteLUT[7816] = 16'h82aa;
RsqrteLUT[7817] = 16'h82a5;
RsqrteLUT[7818] = 16'h82a1;
RsqrteLUT[7819] = 16'h829c;
RsqrteLUT[7820] = 16'h8298;
RsqrteLUT[7821] = 16'h8294;
RsqrteLUT[7822] = 16'h828f;
RsqrteLUT[7823] = 16'h828b;
RsqrteLUT[7824] = 16'h8287;
RsqrteLUT[7825] = 16'h8283;
RsqrteLUT[7826] = 16'h827f;
RsqrteLUT[7827] = 16'h827b;
RsqrteLUT[7828] = 16'h8278;
RsqrteLUT[7829] = 16'h8274;
RsqrteLUT[7830] = 16'h8270;
RsqrteLUT[7831] = 16'h826d;
RsqrteLUT[7832] = 16'h8269;
RsqrteLUT[7833] = 16'h8266;
RsqrteLUT[7834] = 16'h8262;
RsqrteLUT[7835] = 16'h825f;
RsqrteLUT[7836] = 16'h825b;
RsqrteLUT[7837] = 16'h8258;
RsqrteLUT[7838] = 16'h8255;
RsqrteLUT[7839] = 16'h8252;
RsqrteLUT[7840] = 16'h824f;
RsqrteLUT[7841] = 16'h824c;
RsqrteLUT[7842] = 16'h8249;
RsqrteLUT[7843] = 16'h8246;
RsqrteLUT[7844] = 16'h8243;
RsqrteLUT[7845] = 16'h8240;
RsqrteLUT[7846] = 16'h823d;
RsqrteLUT[7847] = 16'h823a;
RsqrteLUT[7848] = 16'h8238;
RsqrteLUT[7849] = 16'h8235;
RsqrteLUT[7850] = 16'h8232;
RsqrteLUT[7851] = 16'h822f;
RsqrteLUT[7852] = 16'h822d;
RsqrteLUT[7853] = 16'h822a;
RsqrteLUT[7854] = 16'h8228;
RsqrteLUT[7855] = 16'h8225;
RsqrteLUT[7856] = 16'h8223;
RsqrteLUT[7857] = 16'h8220;
RsqrteLUT[7858] = 16'h821e;
RsqrteLUT[7859] = 16'h821c;
RsqrteLUT[7860] = 16'h8219;
RsqrteLUT[7861] = 16'h8217;
RsqrteLUT[7862] = 16'h8215;
RsqrteLUT[7863] = 16'h8213;
RsqrteLUT[7864] = 16'h8210;
RsqrteLUT[7865] = 16'h820e;
RsqrteLUT[7866] = 16'h820c;
RsqrteLUT[7867] = 16'h820a;
RsqrteLUT[7868] = 16'h8208;
RsqrteLUT[7869] = 16'h8206;
RsqrteLUT[7870] = 16'h8204;
RsqrteLUT[7871] = 16'h8202;
RsqrteLUT[7872] = 16'h8200;
RsqrteLUT[7873] = 16'h81f8;
RsqrteLUT[7874] = 16'h81f0;
RsqrteLUT[7875] = 16'h81e8;
RsqrteLUT[7876] = 16'h81e1;
RsqrteLUT[7877] = 16'h81da;
RsqrteLUT[7878] = 16'h81d3;
RsqrteLUT[7879] = 16'h81cc;
RsqrteLUT[7880] = 16'h81c5;
RsqrteLUT[7881] = 16'h81be;
RsqrteLUT[7882] = 16'h81b8;
RsqrteLUT[7883] = 16'h81b1;
RsqrteLUT[7884] = 16'h81ab;
RsqrteLUT[7885] = 16'h81a5;
RsqrteLUT[7886] = 16'h819f;
RsqrteLUT[7887] = 16'h8199;
RsqrteLUT[7888] = 16'h8193;
RsqrteLUT[7889] = 16'h818e;
RsqrteLUT[7890] = 16'h8188;
RsqrteLUT[7891] = 16'h8183;
RsqrteLUT[7892] = 16'h817d;
RsqrteLUT[7893] = 16'h8178;
RsqrteLUT[7894] = 16'h8173;
RsqrteLUT[7895] = 16'h816e;
RsqrteLUT[7896] = 16'h8169;
RsqrteLUT[7897] = 16'h8164;
RsqrteLUT[7898] = 16'h815f;
RsqrteLUT[7899] = 16'h815a;
RsqrteLUT[7900] = 16'h8156;
RsqrteLUT[7901] = 16'h8151;
RsqrteLUT[7902] = 16'h814c;
RsqrteLUT[7903] = 16'h8148;
RsqrteLUT[7904] = 16'h8144;
RsqrteLUT[7905] = 16'h813f;
RsqrteLUT[7906] = 16'h813b;
RsqrteLUT[7907] = 16'h8137;
RsqrteLUT[7908] = 16'h8133;
RsqrteLUT[7909] = 16'h812f;
RsqrteLUT[7910] = 16'h812b;
RsqrteLUT[7911] = 16'h8127;
RsqrteLUT[7912] = 16'h8123;
RsqrteLUT[7913] = 16'h811f;
RsqrteLUT[7914] = 16'h811b;
RsqrteLUT[7915] = 16'h8117;
RsqrteLUT[7916] = 16'h8114;
RsqrteLUT[7917] = 16'h8110;
RsqrteLUT[7918] = 16'h810d;
RsqrteLUT[7919] = 16'h8109;
RsqrteLUT[7920] = 16'h8106;
RsqrteLUT[7921] = 16'h8102;
RsqrteLUT[7922] = 16'h80ff;
RsqrteLUT[7923] = 16'h80fb;
RsqrteLUT[7924] = 16'h80f8;
RsqrteLUT[7925] = 16'h80f5;
RsqrteLUT[7926] = 16'h80f2;
RsqrteLUT[7927] = 16'h80ee;
RsqrteLUT[7928] = 16'h80eb;
RsqrteLUT[7929] = 16'h80e8;
RsqrteLUT[7930] = 16'h80e5;
RsqrteLUT[7931] = 16'h80e2;
RsqrteLUT[7932] = 16'h80df;
RsqrteLUT[7933] = 16'h80dc;
RsqrteLUT[7934] = 16'h80d9;
RsqrteLUT[7935] = 16'h80d6;
RsqrteLUT[7936] = 16'h80d4;
RsqrteLUT[7937] = 16'h80ce;
RsqrteLUT[7938] = 16'h80c9;
RsqrteLUT[7939] = 16'h80c3;
RsqrteLUT[7940] = 16'h80be;
RsqrteLUT[7941] = 16'h80b9;
RsqrteLUT[7942] = 16'h80b4;
RsqrteLUT[7943] = 16'h80af;
RsqrteLUT[7944] = 16'h80aa;
RsqrteLUT[7945] = 16'h80a5;
RsqrteLUT[7946] = 16'h80a1;
RsqrteLUT[7947] = 16'h809c;
RsqrteLUT[7948] = 16'h8098;
RsqrteLUT[7949] = 16'h8094;
RsqrteLUT[7950] = 16'h808f;
RsqrteLUT[7951] = 16'h808b;
RsqrteLUT[7952] = 16'h8087;
RsqrteLUT[7953] = 16'h8083;
RsqrteLUT[7954] = 16'h807f;
RsqrteLUT[7955] = 16'h807b;
RsqrteLUT[7956] = 16'h8078;
RsqrteLUT[7957] = 16'h8074;
RsqrteLUT[7958] = 16'h8070;
RsqrteLUT[7959] = 16'h806d;
RsqrteLUT[7960] = 16'h8069;
RsqrteLUT[7961] = 16'h8066;
RsqrteLUT[7962] = 16'h8062;
RsqrteLUT[7963] = 16'h805f;
RsqrteLUT[7964] = 16'h805b;
RsqrteLUT[7965] = 16'h8058;
RsqrteLUT[7966] = 16'h8055;
RsqrteLUT[7967] = 16'h8052;
RsqrteLUT[7968] = 16'h804f;
RsqrteLUT[7969] = 16'h804c;
RsqrteLUT[7970] = 16'h8049;
RsqrteLUT[7971] = 16'h8046;
RsqrteLUT[7972] = 16'h8043;
RsqrteLUT[7973] = 16'h8040;
RsqrteLUT[7974] = 16'h803d;
RsqrteLUT[7975] = 16'h803a;
RsqrteLUT[7976] = 16'h8038;
RsqrteLUT[7977] = 16'h8035;
RsqrteLUT[7978] = 16'h8032;
RsqrteLUT[7979] = 16'h802f;
RsqrteLUT[7980] = 16'h802d;
RsqrteLUT[7981] = 16'h802a;
RsqrteLUT[7982] = 16'h8028;
RsqrteLUT[7983] = 16'h8025;
RsqrteLUT[7984] = 16'h8023;
RsqrteLUT[7985] = 16'h8020;
RsqrteLUT[7986] = 16'h801e;
RsqrteLUT[7987] = 16'h801c;
RsqrteLUT[7988] = 16'h8019;
RsqrteLUT[7989] = 16'h8017;
RsqrteLUT[7990] = 16'h8015;
RsqrteLUT[7991] = 16'h8013;
RsqrteLUT[7992] = 16'h8010;
RsqrteLUT[7993] = 16'h800e;
RsqrteLUT[7994] = 16'h800c;
RsqrteLUT[7995] = 16'h800a;
RsqrteLUT[7996] = 16'h8008;
RsqrteLUT[7997] = 16'h8006;
RsqrteLUT[7998] = 16'h8004;
RsqrteLUT[7999] = 16'h8002;
RsqrteLUT[8000] = 16'h8000;
RsqrteLUT[8001] = 16'h7ff8;
RsqrteLUT[8002] = 16'h7ff0;
RsqrteLUT[8003] = 16'h7fe8;
RsqrteLUT[8004] = 16'h7fe1;
RsqrteLUT[8005] = 16'h7fda;
RsqrteLUT[8006] = 16'h7fd3;
RsqrteLUT[8007] = 16'h7fcc;
RsqrteLUT[8008] = 16'h7fc5;
RsqrteLUT[8009] = 16'h7fbe;
RsqrteLUT[8010] = 16'h7fb8;
RsqrteLUT[8011] = 16'h7fb1;
RsqrteLUT[8012] = 16'h7fab;
RsqrteLUT[8013] = 16'h7fa5;
RsqrteLUT[8014] = 16'h7f9f;
RsqrteLUT[8015] = 16'h7f99;
RsqrteLUT[8016] = 16'h7f93;
RsqrteLUT[8017] = 16'h7f8e;
RsqrteLUT[8018] = 16'h7f88;
RsqrteLUT[8019] = 16'h7f83;
RsqrteLUT[8020] = 16'h7f7d;
RsqrteLUT[8021] = 16'h7f78;
RsqrteLUT[8022] = 16'h7f73;
RsqrteLUT[8023] = 16'h7f6e;
RsqrteLUT[8024] = 16'h7f69;
RsqrteLUT[8025] = 16'h7f64;
RsqrteLUT[8026] = 16'h7f5f;
RsqrteLUT[8027] = 16'h7f5a;
RsqrteLUT[8028] = 16'h7f56;
RsqrteLUT[8029] = 16'h7f51;
RsqrteLUT[8030] = 16'h7f4c;
RsqrteLUT[8031] = 16'h7f48;
RsqrteLUT[8032] = 16'h7f44;
RsqrteLUT[8033] = 16'h7f3f;
RsqrteLUT[8034] = 16'h7f3b;
RsqrteLUT[8035] = 16'h7f37;
RsqrteLUT[8036] = 16'h7f33;
RsqrteLUT[8037] = 16'h7f2f;
RsqrteLUT[8038] = 16'h7f2b;
RsqrteLUT[8039] = 16'h7f27;
RsqrteLUT[8040] = 16'h7f23;
RsqrteLUT[8041] = 16'h7f1f;
RsqrteLUT[8042] = 16'h7f1b;
RsqrteLUT[8043] = 16'h7f17;
RsqrteLUT[8044] = 16'h7f14;
RsqrteLUT[8045] = 16'h7f10;
RsqrteLUT[8046] = 16'h7f0d;
RsqrteLUT[8047] = 16'h7f09;
RsqrteLUT[8048] = 16'h7f06;
RsqrteLUT[8049] = 16'h7f02;
RsqrteLUT[8050] = 16'h7eff;
RsqrteLUT[8051] = 16'h7efb;
RsqrteLUT[8052] = 16'h7ef8;
RsqrteLUT[8053] = 16'h7ef5;
RsqrteLUT[8054] = 16'h7ef2;
RsqrteLUT[8055] = 16'h7eee;
RsqrteLUT[8056] = 16'h7eeb;
RsqrteLUT[8057] = 16'h7ee8;
RsqrteLUT[8058] = 16'h7ee5;
RsqrteLUT[8059] = 16'h7ee2;
RsqrteLUT[8060] = 16'h7edf;
RsqrteLUT[8061] = 16'h7edc;
RsqrteLUT[8062] = 16'h7ed9;
RsqrteLUT[8063] = 16'h7ed6;
RsqrteLUT[8064] = 16'h7ed4;
RsqrteLUT[8065] = 16'h7ece;
RsqrteLUT[8066] = 16'h7ec9;
RsqrteLUT[8067] = 16'h7ec3;
RsqrteLUT[8068] = 16'h7ebe;
RsqrteLUT[8069] = 16'h7eb9;
RsqrteLUT[8070] = 16'h7eb4;
RsqrteLUT[8071] = 16'h7eaf;
RsqrteLUT[8072] = 16'h7eaa;
RsqrteLUT[8073] = 16'h7ea5;
RsqrteLUT[8074] = 16'h7ea1;
RsqrteLUT[8075] = 16'h7e9c;
RsqrteLUT[8076] = 16'h7e98;
RsqrteLUT[8077] = 16'h7e94;
RsqrteLUT[8078] = 16'h7e8f;
RsqrteLUT[8079] = 16'h7e8b;
RsqrteLUT[8080] = 16'h7e87;
RsqrteLUT[8081] = 16'h7e83;
RsqrteLUT[8082] = 16'h7e7f;
RsqrteLUT[8083] = 16'h7e7b;
RsqrteLUT[8084] = 16'h7e78;
RsqrteLUT[8085] = 16'h7e74;
RsqrteLUT[8086] = 16'h7e70;
RsqrteLUT[8087] = 16'h7e6d;
RsqrteLUT[8088] = 16'h7e69;
RsqrteLUT[8089] = 16'h7e66;
RsqrteLUT[8090] = 16'h7e62;
RsqrteLUT[8091] = 16'h7e5f;
RsqrteLUT[8092] = 16'h7e5b;
RsqrteLUT[8093] = 16'h7e58;
RsqrteLUT[8094] = 16'h7e55;
RsqrteLUT[8095] = 16'h7e52;
RsqrteLUT[8096] = 16'h7e4f;
RsqrteLUT[8097] = 16'h7e4c;
RsqrteLUT[8098] = 16'h7e49;
RsqrteLUT[8099] = 16'h7e46;
RsqrteLUT[8100] = 16'h7e43;
RsqrteLUT[8101] = 16'h7e40;
RsqrteLUT[8102] = 16'h7e3d;
RsqrteLUT[8103] = 16'h7e3a;
RsqrteLUT[8104] = 16'h7e38;
RsqrteLUT[8105] = 16'h7e35;
RsqrteLUT[8106] = 16'h7e32;
RsqrteLUT[8107] = 16'h7e2f;
RsqrteLUT[8108] = 16'h7e2d;
RsqrteLUT[8109] = 16'h7e2a;
RsqrteLUT[8110] = 16'h7e28;
RsqrteLUT[8111] = 16'h7e25;
RsqrteLUT[8112] = 16'h7e23;
RsqrteLUT[8113] = 16'h7e20;
RsqrteLUT[8114] = 16'h7e1e;
RsqrteLUT[8115] = 16'h7e1c;
RsqrteLUT[8116] = 16'h7e19;
RsqrteLUT[8117] = 16'h7e17;
RsqrteLUT[8118] = 16'h7e15;
RsqrteLUT[8119] = 16'h7e13;
RsqrteLUT[8120] = 16'h7e10;
RsqrteLUT[8121] = 16'h7e0e;
RsqrteLUT[8122] = 16'h7e0c;
RsqrteLUT[8123] = 16'h7e0a;
RsqrteLUT[8124] = 16'h7e08;
RsqrteLUT[8125] = 16'h7e06;
RsqrteLUT[8126] = 16'h7e04;
RsqrteLUT[8127] = 16'h7e02;
RsqrteLUT[8128] = 16'h7e00;
RsqrteLUT[8129] = 16'h7df8;
RsqrteLUT[8130] = 16'h7df0;
RsqrteLUT[8131] = 16'h7de8;
RsqrteLUT[8132] = 16'h7de1;
RsqrteLUT[8133] = 16'h7dda;
RsqrteLUT[8134] = 16'h7dd3;
RsqrteLUT[8135] = 16'h7dcc;
RsqrteLUT[8136] = 16'h7dc5;
RsqrteLUT[8137] = 16'h7dbe;
RsqrteLUT[8138] = 16'h7db8;
RsqrteLUT[8139] = 16'h7db1;
RsqrteLUT[8140] = 16'h7dab;
RsqrteLUT[8141] = 16'h7da5;
RsqrteLUT[8142] = 16'h7d9f;
RsqrteLUT[8143] = 16'h7d99;
RsqrteLUT[8144] = 16'h7d93;
RsqrteLUT[8145] = 16'h7d8e;
RsqrteLUT[8146] = 16'h7d88;
RsqrteLUT[8147] = 16'h7d83;
RsqrteLUT[8148] = 16'h7d7d;
RsqrteLUT[8149] = 16'h7d78;
RsqrteLUT[8150] = 16'h7d73;
RsqrteLUT[8151] = 16'h7d6e;
RsqrteLUT[8152] = 16'h7d69;
RsqrteLUT[8153] = 16'h7d64;
RsqrteLUT[8154] = 16'h7d5f;
RsqrteLUT[8155] = 16'h7d5a;
RsqrteLUT[8156] = 16'h7d56;
RsqrteLUT[8157] = 16'h7d51;
RsqrteLUT[8158] = 16'h7d4c;
RsqrteLUT[8159] = 16'h7d48;
RsqrteLUT[8160] = 16'h7d44;
RsqrteLUT[8161] = 16'h7d3f;
RsqrteLUT[8162] = 16'h7d3b;
RsqrteLUT[8163] = 16'h7d37;
RsqrteLUT[8164] = 16'h7d33;
RsqrteLUT[8165] = 16'h7d2f;
RsqrteLUT[8166] = 16'h7d2b;
RsqrteLUT[8167] = 16'h7d27;
RsqrteLUT[8168] = 16'h7d23;
RsqrteLUT[8169] = 16'h7d1f;
RsqrteLUT[8170] = 16'h7d1b;
RsqrteLUT[8171] = 16'h7d17;
RsqrteLUT[8172] = 16'h7d14;
RsqrteLUT[8173] = 16'h7d10;
RsqrteLUT[8174] = 16'h7d0d;
RsqrteLUT[8175] = 16'h7d09;
RsqrteLUT[8176] = 16'h7d06;
RsqrteLUT[8177] = 16'h7d02;
RsqrteLUT[8178] = 16'h7cff;
RsqrteLUT[8179] = 16'h7cfb;
RsqrteLUT[8180] = 16'h7cf8;
RsqrteLUT[8181] = 16'h7cf5;
RsqrteLUT[8182] = 16'h7cf2;
RsqrteLUT[8183] = 16'h7cee;
RsqrteLUT[8184] = 16'h7ceb;
RsqrteLUT[8185] = 16'h7ce8;
RsqrteLUT[8186] = 16'h7ce5;
RsqrteLUT[8187] = 16'h7ce2;
RsqrteLUT[8188] = 16'h7cdf;
RsqrteLUT[8189] = 16'h7cdc;
RsqrteLUT[8190] = 16'h7cd9;
RsqrteLUT[8191] = 16'h7cd6;
end

wire [31:0] a1;
reg [31:0] o1;
reg s1, s2;
F80ToF32 u1 (a, a1);
F32ToF80 u2 (o1, o);

wire [13:0] index = a1[30:17];
reg [13:0] indexr;
reg [16:0] luto;


always @(posedge clk)
	if (ce) indexr <= index;
always @(posedge clk)
	if(ce) s1 <= a1[31];
always @(posedge clk)
if (ce) begin
	s2 <= s1;
	if (indexr < 14'd8129)
		luto <= 17'h7FC0 << 1;
	else if (indexr < 14'd8197)
		luto <= RsqrteLUT2[indexr - 14'd8197] << 1;
	else
		luto <= RsqrteLUT[indexr[12:0]];
end

wire [7:0] exp = luto[16:9];
wire [22:0] man = {luto[8:0],14'd0};
always @*
	if (s2)
		o1 <= {1'b0,`QSQRTNEG};
	else
		o1 = {1'b0,exp,man};

`else
`ifdef RSQRT_SM
// Reciprocal square root estimate using a state machine.

wire [31:0] a1;
reg [31:0] x2, x2yy;
reg [31:0] y, yy;
wire [31:0] y1 = `FRSQRTE_MAGIC - a1[31:1];
reg [31:0] aa0, bb0, aa1, bb1;
wire [31:0] mo0, mo1, x2yy1p5;

reg [3:0] cnt;
reg [2:0] state;
parameter IDLE = 3'd0;
parameter MULP5 = 3'd1;
parameter MULX2YY = 3'd2;
parameter SUB = 3'd3;
parameter RES = 3'd4;

always @(posedge clk)
begin
	if (ld) begin
		state <= MULP5;
		cnt <= 4'd5;
		aa0 <= a1;
		bb0 <= `POINT5;
		aa1 <= y1;
		bb1 <= y1;
		y <= y1;
	end
	case(state)
	IDLE:	;
	MULP5:	
		begin
			cnt <= cnt - 4'd1;
			if (cnt[3]) begin
				cnt <= 4'd5;
				x2 <= mo0;
				yy <= mo1;
				aa0 <= mo0;
				bb0 <= mo1;
				state <= MULX2YY;
			end
		end
	MULX2YY:
		begin
			cnt <= cnt - 4'd1;
			if (cnt[3]) begin
				cnt <= 4'd5;
				x2yy <= mo0;
				aa0 <= `ONEPOINT5;
				bb0 <= mo0;
				state <= SUB;
			end
		end
	SUB:
		begin
			cnt <= cnt - 4'd1;
			if (cnt[3]) begin
				cnt <= 4'd5;
				aa0 <= y;
				bb0 <= x2yy1p5;
				state <= RES;
			end
		end
	RES:
		begin
			cnt <= cnt - 4'd1;
			if (cnt[3]) begin
				state <= IDLE;
			end
		end
	endcase
end

F80ToF32 u0 (a, a1);
fpMulnr #(32) u1 (clk, ce, aa0, bb0, mo0);
fpMulnr #(32) u2 (clk, ce, aa1, bb1, mo1);
fpAddsubnr #(32) u3 (clk, ce, 3'd0, 1'b1, aa0, bb0, x2yy1p5);
F32ToF80 u4 (mo0, o);

`else
// Reciprocal square root estimate using FP hardware.

fpMulnr #(32) u1 (clk, ce, a, `POINT5, x2);
assign y = `FRSQRTE_MAGIC - a[31:1];
fpMulnr #(32) u2 (clk, ce, y, y, yy);
fpMulnr #(32) u3 (clk, ce, x2, yy, x2yy);
fpAddsubnr #(32) u4 (clk, ce, 3'd0, 1'b1, `ONEPOINT5, x2yy, x2yy1p5);
fpMulnr #(32) u5 (clk, ce, y, x2yy1p5, o);

`endif
`endif

endmodule
